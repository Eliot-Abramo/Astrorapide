version https://git-lfs.github.com/spec/v1
oid sha256:bfa06000de02d7cf6e51f3261724c63353d1ad908f17bc1125b5dc38d3d937c2
size 54070
