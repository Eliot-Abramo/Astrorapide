version https://git-lfs.github.com/spec/v1
oid sha256:a3e79335c95d899d0cc91afc2f2c337bb8bd8c055a15baa934112f278e0b91da
size 20964
