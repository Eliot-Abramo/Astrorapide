version https://git-lfs.github.com/spec/v1
oid sha256:375687e42853e59a9b4851e8618df04d93d249118685caca822a499e9de36294
size 4487
