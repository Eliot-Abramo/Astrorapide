version https://git-lfs.github.com/spec/v1
oid sha256:ae5944fb786659eae6dc8f9b69f30fa920e7628b3e314e9747653a21bdf68762
size 13250
