version https://git-lfs.github.com/spec/v1
oid sha256:caf8ee77b5058899609e8f947ca1fe56fac15afafd23936a6f35f7d5ff15f462
size 14667
