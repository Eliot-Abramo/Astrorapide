version https://git-lfs.github.com/spec/v1
oid sha256:34bf051503e6140fb176dd961619593651364c4a33aefd5b708933f1769c0da3
size 2106
