version https://git-lfs.github.com/spec/v1
oid sha256:2f8e810debcc20834e201616e27b4f5fd8b7aed957b02d758eeae693924a6943
size 48277
