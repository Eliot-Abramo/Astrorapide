version https://git-lfs.github.com/spec/v1
oid sha256:e028ec5a66040b250923e1ac84ef7b6f5f596de8e323e6211c177d8237ee6586
size 4491
