version https://git-lfs.github.com/spec/v1
oid sha256:eee76b1fb4a60185ee1eac92ceedefd42d7b409929bdd4989ec8278668672f48
size 2843
