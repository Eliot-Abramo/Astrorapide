version https://git-lfs.github.com/spec/v1
oid sha256:ef80658eb913a1668a556db6c79ad125ff410a2dad0822d1c39b7ff327c0c190
size 2111
