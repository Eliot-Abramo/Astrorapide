version https://git-lfs.github.com/spec/v1
oid sha256:4e3368f3fe8a0fb3718c043f00f14aab87c1a18a68d30c0a11141e53243ea8cf
size 2108
