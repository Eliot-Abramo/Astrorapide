version https://git-lfs.github.com/spec/v1
oid sha256:fdecdf3ddb7df9d906b2e002bda9cdd01961e099bd23ee6fe6ad44d47dc4f275
size 12952
