version https://git-lfs.github.com/spec/v1
oid sha256:64a4d4bb1f3bcc70c71ef2b055f7fe7703c5e4ba3207a459f7b05d6596925769
size 14332
