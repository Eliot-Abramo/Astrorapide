version https://git-lfs.github.com/spec/v1
oid sha256:d525bbc23c5a0fb9cc11d66910fdd586f4231a0961b15a023cbaebe1f23d2c86
size 24472
