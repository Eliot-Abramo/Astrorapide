version https://git-lfs.github.com/spec/v1
oid sha256:fb96dda32c0d213e14575af2149098b8e65b32b1d35d0fa779b16104ecde2c12
size 113822
