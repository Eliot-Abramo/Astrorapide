version https://git-lfs.github.com/spec/v1
oid sha256:ad1dc8d4c7cad55d2d9523016e08851a6878da0d6197e92d5e8916fe5e75741b
size 5313
