version https://git-lfs.github.com/spec/v1
oid sha256:e88e159df91aed3f7f78824cc0edefcaf9905c4fc54c804221c72d8f5a219c6d
size 13373
