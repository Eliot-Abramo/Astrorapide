version https://git-lfs.github.com/spec/v1
oid sha256:44fdb9014a4dac07b68d74bd3543ecb661e38fceb91e59e4d835197c7fbfd928
size 13386
