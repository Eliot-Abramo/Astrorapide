version https://git-lfs.github.com/spec/v1
oid sha256:7f47b57b39b36f3a913078eb9644fe32cb6d5ef55209b352374a840f4b82df9a
size 14336
