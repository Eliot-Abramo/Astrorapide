version https://git-lfs.github.com/spec/v1
oid sha256:fe88e1c4803579373c9292fad7c34ae1c10357c43f0e733759ad90f9abf34bce
size 43958
