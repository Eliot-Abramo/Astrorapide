version https://git-lfs.github.com/spec/v1
oid sha256:6b217a3bfdb2b0478ad7a8562831731d6375d94f41a467c6a4e56dda0a869ef5
size 14535
