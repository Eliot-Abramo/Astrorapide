version https://git-lfs.github.com/spec/v1
oid sha256:0d5d0f117e21bd84960a465aa7bd773737ed78443264825a43859feeb57c4797
size 25584
