version https://git-lfs.github.com/spec/v1
oid sha256:3832f05e90a57d44bf83c03efa193024676edd097204dadd70c4c1299d1f4f39
size 1194
