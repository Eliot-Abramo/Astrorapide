version https://git-lfs.github.com/spec/v1
oid sha256:f97556804cbeb7f04f0843c423708f1683d9e1bdcab52666aa2eed59b5772987
size 43396
