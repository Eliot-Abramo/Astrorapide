version https://git-lfs.github.com/spec/v1
oid sha256:969e5459ae978d1b644aab528ffdae46d7ad05be76c64856f2889b30929dc12e
size 14500
