version https://git-lfs.github.com/spec/v1
oid sha256:16461f45cce055afcda404eba6d18582ec34f6768218141878be72aa334e20da
size 1809
