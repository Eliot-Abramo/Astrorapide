version https://git-lfs.github.com/spec/v1
oid sha256:dd6cb5254867997cdce998e1aa6df8ba70ba87802bd1878489a50c7eb2898733
size 30880
