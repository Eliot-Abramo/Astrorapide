version https://git-lfs.github.com/spec/v1
oid sha256:fc12e7d1f3678139b5ad2bac57c0eb9b00d517a1c48b6707fb26d9a85946d333
size 2826
