version https://git-lfs.github.com/spec/v1
oid sha256:730695a9a9a027cc74c68e22686b635c105e53d61f88764c51463055e34e0f70
size 81212
