version https://git-lfs.github.com/spec/v1
oid sha256:1fc98aff1592f43f6c86bb5a0a21bdd0e8ea733f5bee8694e8a1bf9f7de27f46
size 9977
