version https://git-lfs.github.com/spec/v1
oid sha256:175bdccb506c1836444083ca0553d9955730f7418d9d867a46cf30b26de8df40
size 2836
