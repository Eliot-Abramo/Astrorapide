version https://git-lfs.github.com/spec/v1
oid sha256:c826a50d72f818a5fcafba7ce4f25dd47eb8c120fa7996165f79eec3436f0b30
size 17439
