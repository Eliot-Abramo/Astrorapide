version https://git-lfs.github.com/spec/v1
oid sha256:8009f6102d7f4aaa9de4f0cc8affa7b4a018696b38e760eeb3dfdc1a632a65e9
size 5542
