version https://git-lfs.github.com/spec/v1
oid sha256:936a91a23203f928e943085551dadfcd8954450f7170645625e5ba2781187c59
size 12530
