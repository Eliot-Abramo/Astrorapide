version https://git-lfs.github.com/spec/v1
oid sha256:483e042e50c1bae56c9db1a94db5831583b4242bd9a286800c89bf075a6831cc
size 108589
