version https://git-lfs.github.com/spec/v1
oid sha256:78ecece06cb8336a9ce83614131726426f9355978ad921b43bd648b6cd4f6bb3
size 54967
