version https://git-lfs.github.com/spec/v1
oid sha256:699f5ba151e4190c4e9f65256fe3957fe8a41f7bf246148066461d2b0a67efd5
size 44499
