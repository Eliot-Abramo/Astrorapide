version https://git-lfs.github.com/spec/v1
oid sha256:1d1382d54d1fa46285853c041f4808c013ffd883a290d3f14357802987442211
size 86285
