version https://git-lfs.github.com/spec/v1
oid sha256:86e03a57bba6a2ec1acc8e8c0e636e5404d5aed663de4b54b7cefc035020cf01
size 10096
