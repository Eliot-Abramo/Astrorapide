version https://git-lfs.github.com/spec/v1
oid sha256:2678ca29b6301f3d253551d173b9482ea9e12ce919c4fcf2bb46f0f929a51772
size 49371
