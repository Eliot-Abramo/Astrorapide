version https://git-lfs.github.com/spec/v1
oid sha256:1861723e7d05359b64c53694408eae110bcb28caee3df84008eb4749c9011bcc
size 43930
