version https://git-lfs.github.com/spec/v1
oid sha256:ed38840813e8a52475302888f6e8e0b3e7610412dd8598b6b6fe9727c626127c
size 18537
