version https://git-lfs.github.com/spec/v1
oid sha256:6aea175b2633af7aab3337b3e2eaaf1debd74f825fd7a6ff0a628494bcb6d7cc
size 25584
