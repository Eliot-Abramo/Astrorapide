version https://git-lfs.github.com/spec/v1
oid sha256:7e03085a316a88026043902143b7e7554494ba1b79fb30cb063412f5e0323279
size 61032
