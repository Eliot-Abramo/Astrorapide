version https://git-lfs.github.com/spec/v1
oid sha256:dfadd41be39c39469c04c64855a78471a05bd5fb838d4196c4e5ae552f51b1fc
size 14528
