version https://git-lfs.github.com/spec/v1
oid sha256:dc9a8e0ac686ed24ac8cb891999c0b9711cbc63d8b442b5f3a42dc53954df178
size 2849
