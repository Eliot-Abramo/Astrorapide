version https://git-lfs.github.com/spec/v1
oid sha256:68b55ec5a813a5c9ed0c6ecbd8bcb34bcba0713f7c7b41bbf6da9b33b9fae58d
size 54893
