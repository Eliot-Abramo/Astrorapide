version https://git-lfs.github.com/spec/v1
oid sha256:eca3c5aa2b320d57e28c2b1da9488354ee79b2f523a1bc43c32693727ea70d32
size 2054
