version https://git-lfs.github.com/spec/v1
oid sha256:100b56bbcfb4a00c79b18b48d07b1a53fae8953343d391836a5ec15d0d01e682
size 13470
