version https://git-lfs.github.com/spec/v1
oid sha256:1d260413a6539804054bed2827682ed7d330bd4d9b73c024766cd9d38602372c
size 2840
