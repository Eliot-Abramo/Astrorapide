version https://git-lfs.github.com/spec/v1
oid sha256:04636c32468a6e334038ad74c64fabe0169d3738e6babbbe619aa29a840c4a5a
size 14528
