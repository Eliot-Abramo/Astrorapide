version https://git-lfs.github.com/spec/v1
oid sha256:9c02abaed0d8159a91824efd0b61c9d8da0f22af886980da81edbe440d890251
size 68781
