version https://git-lfs.github.com/spec/v1
oid sha256:658bceadc615410eccad879c1be6b083d4abb5a97dfb5f39b3d13cc3739aed07
size 13183
