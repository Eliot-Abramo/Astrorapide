version https://git-lfs.github.com/spec/v1
oid sha256:8b92c033fe63f5e1c28023b669a0860ccd32867e0166efc983d5bd61899892e8
size 48770
