version https://git-lfs.github.com/spec/v1
oid sha256:ece02ff9794ff40596b78d092084d91e23b5349422d3409629f8790d64b66f5e
size 3654
