version https://git-lfs.github.com/spec/v1
oid sha256:7b200da08de714ebaf5750aa933ee4e47a449c3fb8ec81ff980e19e120d3ef73
size 1809
