version https://git-lfs.github.com/spec/v1
oid sha256:071775b43cb5024602dcd58ad352fdffaeca3ab7cb5d56cf014c7784ead70db2
size 54314
