version https://git-lfs.github.com/spec/v1
oid sha256:a04140e95638c7a4e04fb82e42e5976ed7645680a6abed010f988ef01ad08da1
size 3915
