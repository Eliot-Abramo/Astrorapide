version https://git-lfs.github.com/spec/v1
oid sha256:0fbe6d442ac3d93c35f2019c4d8f486cada5751f379d78572fd1c8df1735dc56
size 75514
