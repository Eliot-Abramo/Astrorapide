version https://git-lfs.github.com/spec/v1
oid sha256:bbbacfbc291e7ce665da6564125e3bd309a542240ef34066ec7b8b92e7c0dc3a
size 93298
