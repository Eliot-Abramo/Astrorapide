version https://git-lfs.github.com/spec/v1
oid sha256:c594eb965854326b3982121d0b3a808cbef869cd124c72af25bee80a3da42f52
size 19678
