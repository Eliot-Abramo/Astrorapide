version https://git-lfs.github.com/spec/v1
oid sha256:63a78cf1bd8a403a39cc137fa5a10d91d8d1207d4f4d6c183e967b215c23267d
size 24470
