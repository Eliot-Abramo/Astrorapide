version https://git-lfs.github.com/spec/v1
oid sha256:ebf7ad4c8f80049c957f84c782b7fdd5cf69f168dc3d817f048db328e2418c3c
size 24470
