version https://git-lfs.github.com/spec/v1
oid sha256:6173dda36bd2c587cc6378c36069e02f8f9f8c07ec4c8326bc7e395aec268143
size 1889
