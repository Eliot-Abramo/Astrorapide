version https://git-lfs.github.com/spec/v1
oid sha256:1c1e088513260de44d90dbff6e3595a9e726f576bf4eab657f84deaa8f3d9554
size 10904
