version https://git-lfs.github.com/spec/v1
oid sha256:054abd35aa7189cf0753a32c4a1e5f63dbfb9ddc38aa01cdfbd6abfb2f0d2b39
size 12482
