version https://git-lfs.github.com/spec/v1
oid sha256:a837b694f6a0bda55997f00e3616dabfefe65a8899f20eacf96954afc68a3272
size 17649
