version https://git-lfs.github.com/spec/v1
oid sha256:8e5553ded307bed9a0354a0052782fd082f835cd120d0e42840a36572d4692f8
size 1180
