version https://git-lfs.github.com/spec/v1
oid sha256:c1c214c4f61fcdf83af0f7783c43d41d7ddea64a9ceb24b2e23d315f43b56528
size 13404
