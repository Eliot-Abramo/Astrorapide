version https://git-lfs.github.com/spec/v1
oid sha256:3b4392cde9c9c17356f07c90c560595e36773b5254b55d4269ecf8a1a5bd13ee
size 113834
