version https://git-lfs.github.com/spec/v1
oid sha256:a1137c34e092d0436801f48c5dcc6cc890fbfa682f7c81a7c2f44e8da17257a1
size 43956
