version https://git-lfs.github.com/spec/v1
oid sha256:bad0ea955de4f636fb0654a666c8d00a8e0852d71dc0d2d1f5d4312d192b8707
size 2086
