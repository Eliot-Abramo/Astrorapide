version https://git-lfs.github.com/spec/v1
oid sha256:8cfb8ce7a41e1d0d664410933d5affcdd012f20e1c532f9f64788bde754ffb4c
size 2116
