version https://git-lfs.github.com/spec/v1
oid sha256:5af1be38a4a98dab8dc94766bb0fe511992a8019b5574794b8a1d439a2fc51c7
size 2107
