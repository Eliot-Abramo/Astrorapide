version https://git-lfs.github.com/spec/v1
oid sha256:73ec40844c15d42a75e11c0ccd45f42663f704891499ffbd0debe6732fdd4ca8
size 43934
