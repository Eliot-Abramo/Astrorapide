version https://git-lfs.github.com/spec/v1
oid sha256:85280e0bd5faad778b5694203b93e9582845f2da08de3f45332b86c8c975f2f1
size 1807
