version https://git-lfs.github.com/spec/v1
oid sha256:ba21a654ed2273a99c3bc703baf0dc1fc48ae55bd61498fe0f7d5929f8102e40
size 51777
