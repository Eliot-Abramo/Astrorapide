version https://git-lfs.github.com/spec/v1
oid sha256:0b5337c7b221e306e536730f5cc3a4b847cd2f78ab6ae32f6dc219233b94cbf1
size 13558
