version https://git-lfs.github.com/spec/v1
oid sha256:a1dd5dcf8e5c16106a43b3e1de04f5c872e3c810efbd0e52306f3492fad5c67a
size 5313
