version https://git-lfs.github.com/spec/v1
oid sha256:36e184865b7905e06677cd1b08e397ae3fd25d4713a86ef7d5379310f18f31aa
size 2819
