version https://git-lfs.github.com/spec/v1
oid sha256:912450a25fed57162443675459403c21e31a3e9f62f23b88d62279ab044351d5
size 17649
