version https://git-lfs.github.com/spec/v1
oid sha256:243ef902742055c967cb867181ace16d410b60704bada05731958eeff227737a
size 38990
