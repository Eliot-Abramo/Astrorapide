version https://git-lfs.github.com/spec/v1
oid sha256:df1a3ca2765b408081f96457675b1bed074c0f615f4c811918c75d32235e2df6
size 2112
