version https://git-lfs.github.com/spec/v1
oid sha256:b2a55ae3b9a3e4f12b9f03c9313143a76b9baa1fb123b8c1260ff1333ef6be4d
size 2415
