version https://git-lfs.github.com/spec/v1
oid sha256:bb7daa5abb76e936e8925fae8f5b29c1c50047a8e8a44553a5faa53248275769
size 2108
