version https://git-lfs.github.com/spec/v1
oid sha256:5e523a0d4a34ab33a2a5c7f900a7b55f3ea17a4f41388ff6bca2b30cafda7414
size 7232
