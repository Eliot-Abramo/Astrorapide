version https://git-lfs.github.com/spec/v1
oid sha256:d4f1547dd5006adb5be19803da0d9b9ea92fd5335d213275d239345b6cc88fc7
size 54848
