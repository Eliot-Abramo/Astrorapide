version https://git-lfs.github.com/spec/v1
oid sha256:dc34bc1d78d9abf1bab1f99b16bafa759147fcb7c113d09a671f0009dce6c4d5
size 20964
