version https://git-lfs.github.com/spec/v1
oid sha256:20ee4fa8466be2e92e2a623cfd59b4aafae0a35c7111dd50ac28b75efe6eebeb
size 42038
