version https://git-lfs.github.com/spec/v1
oid sha256:2d9177ca04fb38f83f7daa59b52e17529d11bead364a0b441b98a2ed53881e02
size 13174
