version https://git-lfs.github.com/spec/v1
oid sha256:7f81a3477b39b6d7e0183fc2b6fd871b5ac47bf1d9dc79a31e04d18668f72b6d
size 19575
