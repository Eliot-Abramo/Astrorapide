version https://git-lfs.github.com/spec/v1
oid sha256:0dcc8efef8a239d152ec42a61292533b15956efca6a180f92809171be4a5d975
size 54941
