version https://git-lfs.github.com/spec/v1
oid sha256:c1e395d9d71e6a330c36abb1e2111ba7b0c27911583bc4c1f60bd18d1d741519
size 43932
