version https://git-lfs.github.com/spec/v1
oid sha256:4b27daf7b7a6b3d2e31b91045efef28c52100625db33418218fe594e73441c05
size 5486
