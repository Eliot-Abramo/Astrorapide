version https://git-lfs.github.com/spec/v1
oid sha256:716ac8815032092738293cffddd2049d442e6d23785db8a4b0ce2f8e8ae5b209
size 19503
