version https://git-lfs.github.com/spec/v1
oid sha256:8a10aeee3e3ef6469a25c5c9f5653dea97c2dd24a786b81452123c5ec30730a6
size 5948
