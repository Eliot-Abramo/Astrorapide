version https://git-lfs.github.com/spec/v1
oid sha256:7318200c0beea1d17b26f52a63a562b05a5430a45a2040ee7e7cc0dabbbfb256
size 9980
