version https://git-lfs.github.com/spec/v1
oid sha256:cb7ba1fc1f56bb32092fb2d48e058e2003864f11457542198dc54d5283d6f36c
size 50837
