version https://git-lfs.github.com/spec/v1
oid sha256:fc5fce82e3ebb9e1cfe1eb7adceb6751aa58343dde85b2296d4b59d3caa7cc5e
size 20970
