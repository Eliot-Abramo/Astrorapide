version https://git-lfs.github.com/spec/v1
oid sha256:81bd5cee29b9f6e32283c7a69c01ba641f3b169e73040bfbcff03c4d6bf02de3
size 13190
