version https://git-lfs.github.com/spec/v1
oid sha256:3bdb33b76b47b56a486f56989c02bf7d534ca40709900d0385108b552914ad6b
size 9981
