version https://git-lfs.github.com/spec/v1
oid sha256:2764579c2aa9934908bc56f1d031436aa59affabef19fc3d831d09fe7fb9e027
size 9978
