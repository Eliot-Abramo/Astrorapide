version https://git-lfs.github.com/spec/v1
oid sha256:19f2c7818a3e6a82b86b537cba190ff11ec3813c13ec85b9d3572364e65bddc8
size 44501
