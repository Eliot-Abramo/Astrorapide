version https://git-lfs.github.com/spec/v1
oid sha256:a94ed38d404535c3dc420ed5543b68a6cb0144d6cd5466d16c1b30bda3699fe3
size 5324
