version https://git-lfs.github.com/spec/v1
oid sha256:f8d00277f82146feff91a11ad2175afd34d3e2069423d4fc8eef0cd38fe42907
size 2412
