version https://git-lfs.github.com/spec/v1
oid sha256:34e94aa6243abbae9315c1e35e3dfdd22f1c3f167a0b5aaa36705789ed9bdf0e
size 5257
