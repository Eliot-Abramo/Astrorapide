version https://git-lfs.github.com/spec/v1
oid sha256:36a0dd6fb46a8ecedc04f29e8d5b2f85805ba5a353eeb3ef6baf334d404ca6b3
size 1871
