version https://git-lfs.github.com/spec/v1
oid sha256:1115abad56ac010f4a48800019a57d33fd1f7aba47397f4a25d1efeb8b6b6077
size 14331
