version https://git-lfs.github.com/spec/v1
oid sha256:512cdbfd48f2f8cc75064e6235b63533633b7a154fe4d92e9ef00a16bea0fb57
size 3659
