version https://git-lfs.github.com/spec/v1
oid sha256:9f66768e7e83a9db86f797274a5cf23beb172bd65f7c80e3ee2ffb0f968ce0d9
size 18135
