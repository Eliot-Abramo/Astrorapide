version https://git-lfs.github.com/spec/v1
oid sha256:6ff81279ee7f468ee63ae550fa1e30e62816b0ac90e89d8564c8cf56be739bef
size 100201
