version https://git-lfs.github.com/spec/v1
oid sha256:faa18038909d38905ecc58471791bd35067c5181dfc060d7611cbd2d20ba2a87
size 13431
