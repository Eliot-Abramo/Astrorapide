version https://git-lfs.github.com/spec/v1
oid sha256:25c81d61a39cef229239ea04b625bb63f74509ad2396237f0b202c7404f3568b
size 5313
