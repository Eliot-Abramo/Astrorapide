version https://git-lfs.github.com/spec/v1
oid sha256:442bce7336fbe9f2bc1199bb08f2dc5b68c344e2ae3e59f60ca31418cc81cb8b
size 14659
