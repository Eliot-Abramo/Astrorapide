version https://git-lfs.github.com/spec/v1
oid sha256:2891e6d05ae2297210ee2fee3f0b1d0c9be602f7b6a207902ab2343262f0e076
size 12938
