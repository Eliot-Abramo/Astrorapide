version https://git-lfs.github.com/spec/v1
oid sha256:fa73ac10fe95ce6978c5ccd08b3d312773a936776db55ed9ff78d0c64f4ec5a7
size 13393
