version https://git-lfs.github.com/spec/v1
oid sha256:0447e15e4d0994fb61529c5b68d14d7caad40b887432a1d9c1729633049aee5b
size 5313
