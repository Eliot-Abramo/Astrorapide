version https://git-lfs.github.com/spec/v1
oid sha256:e5c35c47eb7a648faafc2df59d85ebac608efe8c3ea1ec770a2a44d87da7dc04
size 76095
