version https://git-lfs.github.com/spec/v1
oid sha256:2679c696ac324fdb9e8ede227f20de4fdd3d2c3b912d0837c72e3190d4548ece
size 3277
