version https://git-lfs.github.com/spec/v1
oid sha256:6e251f87d7dbbda2ae60e01110b776679e0f91c36af1ee891b87e72b7cf27369
size 13404
