version https://git-lfs.github.com/spec/v1
oid sha256:5568a0b6e9f17b81b8679c77b3d8e03cb389ee0b020ddc5ddc313ad329f3a81c
size 37766
