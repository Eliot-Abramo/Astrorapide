version https://git-lfs.github.com/spec/v1
oid sha256:1b5e6bc029efff9cabe9f17defedecd16da7f58bbf7a6b4df8c08251379d2d76
size 2843
