version https://git-lfs.github.com/spec/v1
oid sha256:0eb19c6ea57f8a57cc4279e0ef75b1bdd6486cd65528f1813e85a364df6c16e0
size 274952
