version https://git-lfs.github.com/spec/v1
oid sha256:06cd4def8616a098cae99288ca2db18e6f03a9bb27be3b4b2e2e8193dc435497
size 5475
