version https://git-lfs.github.com/spec/v1
oid sha256:9de135c6b9851e93a57eba0895be3839d215e0e515d0e3924463f5543be3f17c
size 49814
