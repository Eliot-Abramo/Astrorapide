version https://git-lfs.github.com/spec/v1
oid sha256:931085027a7d44fea4de0edd33c34316d966cb5770cc7bc77f2b559f26aa4754
size 18713
