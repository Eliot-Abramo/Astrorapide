version https://git-lfs.github.com/spec/v1
oid sha256:76ce58b684bb5d863dfce5c90b99e3dad2d4bf243c568dcc6b1ecb414842a9f0
size 2093
