version https://git-lfs.github.com/spec/v1
oid sha256:5ab253f20e3495f4da0c3fbed283b7f9c350cfdc7a54631cbb4106cf59f2f3e0
size 122987
