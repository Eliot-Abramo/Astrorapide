version https://git-lfs.github.com/spec/v1
oid sha256:0005635726006ca019f93144e347ba46801e9b0e61eec3db91400c0b0e8ef36b
size 12508
