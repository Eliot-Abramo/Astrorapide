version https://git-lfs.github.com/spec/v1
oid sha256:937dde9d9638ac3961710a58d693570c9c0ac2731b19b71b02a49a865209974d
size 2844
