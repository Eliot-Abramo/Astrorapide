version https://git-lfs.github.com/spec/v1
oid sha256:fb85c1084a38ed5b8a44bb9ef8aa789995f941a7b3d7c555a794483f537681b9
size 86303
