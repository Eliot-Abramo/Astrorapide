version https://git-lfs.github.com/spec/v1
oid sha256:206291164a2ac887e7308bb05efff4da864cb8df4fc3ffbf7d00f9288d4dd32b
size 54961
