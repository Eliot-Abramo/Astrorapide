version https://git-lfs.github.com/spec/v1
oid sha256:c160ca5735a78e248b78371ab30a7dc6724bf5ae335b6e8b86e2e5097f216aab
size 5531
