version https://git-lfs.github.com/spec/v1
oid sha256:bef1c70ce427bacfbb1280e1d3e475ddf6623c53d4ef889da069ab2014a7f627
size 111068
