version https://git-lfs.github.com/spec/v1
oid sha256:8a64111a21bb11991f7196a619968c3197569e307582e7825ef189ef6daca399
size 44646
