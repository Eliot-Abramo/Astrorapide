version https://git-lfs.github.com/spec/v1
oid sha256:f8b87da897131b4528ff8546cbca5d707b1a7392c2ab790228d9b242b7725dd8
size 66103
