version https://git-lfs.github.com/spec/v1
oid sha256:d8faa3a15a01f2bbc41327fbbb26e2dac399f4596f77b644b95d22ee7078a473
size 101513
