version https://git-lfs.github.com/spec/v1
oid sha256:51d4401c68c5dfe39dfcb4599d6813616aba272f31b56cb01b2f002b8c415938
size 54179
