version https://git-lfs.github.com/spec/v1
oid sha256:6a54d5ed3ca5b1d4509db58a3461f66f83a1c8018a973d4c458c253f8a5d3d8e
size 20973
