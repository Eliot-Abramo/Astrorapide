version https://git-lfs.github.com/spec/v1
oid sha256:3835063d8140c819c298974fa0722bc07a798cff380f78f5c7c83a8c0d5226f5
size 3659
