version https://git-lfs.github.com/spec/v1
oid sha256:c392e6ce0a0f0c949118e6359e7f908e3733f514df2cb71504bbd76d27a25cc6
size 54189
