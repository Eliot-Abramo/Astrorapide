version https://git-lfs.github.com/spec/v1
oid sha256:bbc28580d45cefddf969cbd87a5e89e0174478b633b229ec8ed8be1aa2df95bd
size 2068
