version https://git-lfs.github.com/spec/v1
oid sha256:406ca277e6653b3c1a83f722f102c77f279b8e5bcd8431fa52ac77ee51664fc3
size 80562
