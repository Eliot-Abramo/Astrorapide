version https://git-lfs.github.com/spec/v1
oid sha256:9fa576378896a2636b7c18a44025a666f29cd30e69ebc2cf7c16d98fb5fc35d4
size 56362
