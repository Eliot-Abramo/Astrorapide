version https://git-lfs.github.com/spec/v1
oid sha256:fa165736ddee9d8d82ed81d0db17862828e2ddc4fa307f7d6de58372d27ba185
size 141307
