version https://git-lfs.github.com/spec/v1
oid sha256:84de36677e2c805d3a39c4430948a1e6f6d4655ea357d58c621e6456457197d4
size 3989
