version https://git-lfs.github.com/spec/v1
oid sha256:4e2f00b3aa8614e60b049465af41a593c9852a57695828ca50a7f31f8f74f472
size 38319
