version https://git-lfs.github.com/spec/v1
oid sha256:28be751663255816c10b77591540206d11b225fb854626cf8dd4e05f16d86605
size 54286
