version https://git-lfs.github.com/spec/v1
oid sha256:5d1f1c1718a3893e0f6a02d90db1b94e325aa15cb8d5b4b8f0c9098e23996a7d
size 3107
