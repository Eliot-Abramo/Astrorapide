version https://git-lfs.github.com/spec/v1
oid sha256:d8a933577a292c53bf9d9114f363766813d3424601aa79114121ccf670b72abe
size 48695
