version https://git-lfs.github.com/spec/v1
oid sha256:9326ae4551381ccddca140534c54b7463afb52384f79ba5df73f80bee4044d55
size 1805
