version https://git-lfs.github.com/spec/v1
oid sha256:41e89ade31ba62ff740bd85b51bcb4740470784d4c9c6f57c444b93f226a8e3d
size 2271
