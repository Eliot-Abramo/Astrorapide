version https://git-lfs.github.com/spec/v1
oid sha256:eb9fad0f46e4baf450f8e5a5a632f5a204a78db8b0e8e2ee60405eb64a27e61f
size 2093
