version https://git-lfs.github.com/spec/v1
oid sha256:9684eec97ae3394cf8b0fc80bb515a93439614bb24810259618e854cf093ff76
size 13467
