version https://git-lfs.github.com/spec/v1
oid sha256:b2e44b111486b5ac4d0252e1b2cfb1932457a850502dee738350378d72c7dfe4
size 2847
