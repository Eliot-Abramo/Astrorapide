version https://git-lfs.github.com/spec/v1
oid sha256:bea89a32f49722576f966573e4c75484886089662d34bed78e486d6254ab371f
size 40111
