version https://git-lfs.github.com/spec/v1
oid sha256:43589d70e8d718fdad1e8179f3034c0c25d141eb547e79ddd085eb782c18fe59
size 43396
