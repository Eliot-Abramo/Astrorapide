version https://git-lfs.github.com/spec/v1
oid sha256:57a08ac7b984cf34a06e2d805ffe5897aef0d99a4c6a36bed817c85a037a3683
size 2840
