version https://git-lfs.github.com/spec/v1
oid sha256:57272d1e63c357c426d22f9fe19bcd8c9cf25488ed07c633e287f80abccac17f
size 18004
