version https://git-lfs.github.com/spec/v1
oid sha256:cd64385d9804b42b587ae40adfecd65d161574b97a26a3bf272071332e09b9c8
size 5257
