version https://git-lfs.github.com/spec/v1
oid sha256:b622a98d8fbee15503261da1c4ea35f260f5c5157efdb602621d693dc8ae28c1
size 2835
