version https://git-lfs.github.com/spec/v1
oid sha256:11471db8bd183ef9541f24c52fa2a08aa426050396d40629575e6defaa8b51ba
size 13379
