version https://git-lfs.github.com/spec/v1
oid sha256:a5da54f0464648338649520458c6aab95a5505245b9dbeb991435554d51c043c
size 1996
