version https://git-lfs.github.com/spec/v1
oid sha256:cd6e6b3789ac77182971bf116721a7f8e9b6177d2956643cc2244b280961a8d7
size 50103
