version https://git-lfs.github.com/spec/v1
oid sha256:ee2490c26e41d7133c315f9869de192222a8a55476a6b853d0333cbcc649631c
size 54130
