version https://git-lfs.github.com/spec/v1
oid sha256:e805afa08a8edfc04c98c9f0923d68d3fc5c2111a6ba98e6d43b3564df87b6c2
size 13407
