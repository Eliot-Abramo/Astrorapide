version https://git-lfs.github.com/spec/v1
oid sha256:48539e3bbb9ee68c5a4fdb30e5c1d309997b7b162312f5d3b05e052f41d4f3c4
size 19752
