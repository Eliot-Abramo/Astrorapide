version https://git-lfs.github.com/spec/v1
oid sha256:1089af593bdaaffd6087919302b6c0981c26f33d4c0ee9502609779ec7c2dde0
size 13387
