version https://git-lfs.github.com/spec/v1
oid sha256:c4952ab756c90dc9af3515baccdc6189e56906f919c89acb6769614fb8df8673
size 14415
