version https://git-lfs.github.com/spec/v1
oid sha256:fb3f9c8d7c36d6c9f5d521737e05487c8b200c8e5c391da8e48332c61dfb726a
size 14664
