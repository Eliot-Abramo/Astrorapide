version https://git-lfs.github.com/spec/v1
oid sha256:c57106fc43e0dc0ee029188ca8078ad9d5431030f7ac9d5b65dc991edef158a3
size 79130
