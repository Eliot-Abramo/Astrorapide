version https://git-lfs.github.com/spec/v1
oid sha256:799ee4f259d5df9f4c38ad87ea102053bb48e725e62827ff5885be8482e32978
size 3105
