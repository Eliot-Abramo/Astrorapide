version https://git-lfs.github.com/spec/v1
oid sha256:4c9d8cdb46014ababd11c7449eb26e2d815f31aa2d50a0814d94747258cf0735
size 43956
