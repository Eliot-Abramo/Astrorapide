version https://git-lfs.github.com/spec/v1
oid sha256:d37941f094fdddf272494ad9cf0ad8d521928a12a2929eb39fe049d5470bcec3
size 54167
