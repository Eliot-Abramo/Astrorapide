version https://git-lfs.github.com/spec/v1
oid sha256:6e0b4de2b664a7deef66381a286ad36ba8f25bcef8971eff1b7fe1508bafd270
size 50923
