version https://git-lfs.github.com/spec/v1
oid sha256:63ba41d3a9389192de0de8e9a6250b2c86fe77acb41c5360f87fd1d878ce1036
size 2426
