version https://git-lfs.github.com/spec/v1
oid sha256:aa28885630f6365296fc4dfa03cff0b2addd21d58531846dcf2af3273929e6f3
size 2108
