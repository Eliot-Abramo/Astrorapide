version https://git-lfs.github.com/spec/v1
oid sha256:aee50dfa85a3d0b283228b30f59dc29f7eb454940a696c9e810d54cefc165e6a
size 1755
