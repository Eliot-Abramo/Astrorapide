version https://git-lfs.github.com/spec/v1
oid sha256:e02dfc3103d8e14fea5269374ced345c0df7ff1b27a35caecb65e2d265ad0808
size 17002
