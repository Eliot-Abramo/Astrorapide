version https://git-lfs.github.com/spec/v1
oid sha256:5b78bf74e77e31f4b090220d67c248ec7dc886b813145492a9a0117a9def30e8
size 1823
