version https://git-lfs.github.com/spec/v1
oid sha256:26417499d1f0704d0353b979ad4ba532cbe999e0faf250f51656150d094f3a38
size 5380
