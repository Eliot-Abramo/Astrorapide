version https://git-lfs.github.com/spec/v1
oid sha256:0e666eab3f2b5ee05b0cf52a93d6cca91ccf10a4f86a914ae01da7599778be46
size 13038
