version https://git-lfs.github.com/spec/v1
oid sha256:ac57e44e4e1ab6997c97e8cea86543c7429802cf58419988f51f3fae49952b19
size 18732
