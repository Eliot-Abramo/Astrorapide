version https://git-lfs.github.com/spec/v1
oid sha256:d49d9b0d6f3a1036dbad6a9951a19e109cd510815c4421bec1e01788c92067a5
size 7284
