version https://git-lfs.github.com/spec/v1
oid sha256:a31e832299627888185773f0bb21149417abc0db68d63c455cc748dec697200d
size 14524
