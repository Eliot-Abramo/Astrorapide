version https://git-lfs.github.com/spec/v1
oid sha256:a829a2f80c7a64f07ba254b9ea52e28c06e85f346e423691feb7d2680a48f19a
size 49489
