version https://git-lfs.github.com/spec/v1
oid sha256:a126ffe0952c9335fa1162daef5586681f545bac9eeb89052d29990c58340d3e
size 2102
