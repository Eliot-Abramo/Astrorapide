version https://git-lfs.github.com/spec/v1
oid sha256:25a9a6b4d999235dd5abb64d4adc4e82d61e55f6833c716d755743d4d95731a1
size 14183
