version https://git-lfs.github.com/spec/v1
oid sha256:59aa783e742118fab3573c225d21ea4416b8549202be2121799e14e870b41ee8
size 9238
