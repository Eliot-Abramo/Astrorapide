version https://git-lfs.github.com/spec/v1
oid sha256:6dfcd0a7204e86ad80f22eb2111a2cbf0bce942bb12db82c06b666a4570d5432
size 3654
