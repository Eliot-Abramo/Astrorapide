version https://git-lfs.github.com/spec/v1
oid sha256:e8316ec5287b64701cba929871215b0967d5639e914c5ceba677dd21614bbb4a
size 5475
