version https://git-lfs.github.com/spec/v1
oid sha256:7a0b9e1d95b8cff89df807472ab8cad7b9b817f40771ef74bf8c255c8f49c175
size 17408
