version https://git-lfs.github.com/spec/v1
oid sha256:de8f397b1793f237bdc58eb0e371e780c7144694359d88d2b2ae42a9d411787f
size 49487
