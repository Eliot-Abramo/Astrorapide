version https://git-lfs.github.com/spec/v1
oid sha256:f300c560e85e238c12aad79240f95a19a861a430bfb9cc5deedc9fdf4eeedadc
size 2102
