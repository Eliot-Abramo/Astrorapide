version https://git-lfs.github.com/spec/v1
oid sha256:efaeab93225b51fc9ce30066059c51bf837156bb40987f8aaec9917700bfc604
size 2068
