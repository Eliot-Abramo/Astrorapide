version https://git-lfs.github.com/spec/v1
oid sha256:61c31af3002ad5b79abc59000639376937e19681f08aedc87cf016f2853edd8f
size 43930
