version https://git-lfs.github.com/spec/v1
oid sha256:dd137d3d55494576d2ecf4fbc46be49a1cdbd2f457d510f12117ba42afe60e65
size 13459
