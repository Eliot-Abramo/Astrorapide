version https://git-lfs.github.com/spec/v1
oid sha256:22f24723bfd6415198d5d59cc8de6e42c8032817650b76aafad00a4f05415d08
size 44495
