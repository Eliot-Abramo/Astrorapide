version https://git-lfs.github.com/spec/v1
oid sha256:5f4b84e013013994e4f09c59052b4ca00ac4a34425614d72e8a921b3bb8493b3
size 25758
