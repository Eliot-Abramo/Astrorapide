version https://git-lfs.github.com/spec/v1
oid sha256:52e6a53a1769246f65e818697d1ea17c045df175e9f9f9f28e928e102f255ba3
size 103344
