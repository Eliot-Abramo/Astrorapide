version https://git-lfs.github.com/spec/v1
oid sha256:256252ef31c6a0ef0cb4f003b94fd213e7437ea53093e35bbf9a1b21a7319e6e
size 2116
