version https://git-lfs.github.com/spec/v1
oid sha256:3947c33b72d46f3b7292f3a4950248ee48d4c2754a273c6e515417ce6528b353
size 2845
