version https://git-lfs.github.com/spec/v1
oid sha256:2d46be0335a1f3e92864ee32406528a351932f15e821ece2c0e6e6bce831d5e0
size 54941
