version https://git-lfs.github.com/spec/v1
oid sha256:60cd7b18d597e89c63aaee1c64e0bd931e41807344a5ab513f2d78423a2bce16
size 2841
