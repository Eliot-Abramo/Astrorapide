version https://git-lfs.github.com/spec/v1
oid sha256:15d9a6d1dfd1254a396e3cd1511e5c15727fafe724ff6e96bda8d80897848dd6
size 13414
