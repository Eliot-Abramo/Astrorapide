version https://git-lfs.github.com/spec/v1
oid sha256:e010161d5b124a54a502238b95a634adc251c0ae26c5c943036f24b4df7ca3d1
size 76095
