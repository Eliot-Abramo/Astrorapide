version https://git-lfs.github.com/spec/v1
oid sha256:f48cc529b5b41695a5f15e2d793b8d4fe3973599d94a8c102fa3202ea8fd3d1f
size 2844
