version https://git-lfs.github.com/spec/v1
oid sha256:7647621008e088be87ab66a87f80125f029626ff7206adfbe4056fb3ec89f1a8
size 13163
