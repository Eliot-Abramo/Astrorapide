version https://git-lfs.github.com/spec/v1
oid sha256:6d33ef4e4c9a3113dc6cfcf7e6e7f4c69f7eddf22900eb45eae38fc88c862476
size 2118
