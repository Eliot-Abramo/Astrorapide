version https://git-lfs.github.com/spec/v1
oid sha256:8f8de1950168867e0ed58da6750fe06db67947f2ad999ffc45e539b9c830c281
size 5321
