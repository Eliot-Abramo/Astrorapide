version https://git-lfs.github.com/spec/v1
oid sha256:8eb6ea23dfb6d4badadc6b0179710c2a49b1ee850cd9cf6ac5ecb2ed973a2a52
size 2100
