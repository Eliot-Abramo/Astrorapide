version https://git-lfs.github.com/spec/v1
oid sha256:dcdc4fbd389cb2e3b0d4b6026e67617925d4742903fa248251592ab6fef0a914
size 76095
