version https://git-lfs.github.com/spec/v1
oid sha256:1ef9618fd56505b6415f78b0bd02d236555afcb17fbdf045d878487864eefacb
size 24286
