version https://git-lfs.github.com/spec/v1
oid sha256:7bb1e623d795d8f62c4929f560b406656ce9e389529f288f9cc797a1e3d1277d
size 21728
