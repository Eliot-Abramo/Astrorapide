version https://git-lfs.github.com/spec/v1
oid sha256:e31c2c8a178194b249a74587e828b2861baf03cb1f087b17abac854be8cf8f85
size 2110
