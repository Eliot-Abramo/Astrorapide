version https://git-lfs.github.com/spec/v1
oid sha256:3a04a2b3bc32ada61dde85c6f07fc6bfc9f192c0a2f60f2d5228e509be273274
size 13398
