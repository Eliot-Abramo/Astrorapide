version https://git-lfs.github.com/spec/v1
oid sha256:4c43f8841887cdd8ee55d9fa5b68121c1003b42968028d2469e4bdeb0c6cf80a
size 3064
