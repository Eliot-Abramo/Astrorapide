version https://git-lfs.github.com/spec/v1
oid sha256:ee06d099cb0c045dcfe399af7dfa5720ec45ff4d212e0c0b83413425c4cf76e8
size 14335
