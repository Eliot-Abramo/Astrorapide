version https://git-lfs.github.com/spec/v1
oid sha256:f89dd70e0e3102c44f2f8f2300944b591898a5dcc20f1649480382a58838776f
size 54286
