version https://git-lfs.github.com/spec/v1
oid sha256:da6b60fc9970c8964fd7c9e01aa82d7b6a7dcc444c22827fc540eca04b32c50d
size 113834
