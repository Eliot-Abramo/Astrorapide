version https://git-lfs.github.com/spec/v1
oid sha256:02f2ca6c2a51f2ef6d08e41a4256f867c87abb121cd06279a72652dc93ed5c08
size 2005
