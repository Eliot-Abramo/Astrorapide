version https://git-lfs.github.com/spec/v1
oid sha256:60c42b9d485ab56a4d95f44d3adea95b0a01608bd9c9097a889141757046b8ff
size 17692
