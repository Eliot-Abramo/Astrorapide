version https://git-lfs.github.com/spec/v1
oid sha256:e5069f9e1ab9dff1db74103ecc7cd8ffe3bb7b7fcdaac84de7037503954de860
size 5257
