version https://git-lfs.github.com/spec/v1
oid sha256:268908682b84e059aebb811fb0f09762d56f6ad2d96d155ec4a31b9692924ed3
size 13166
