version https://git-lfs.github.com/spec/v1
oid sha256:aba18eb31d3ba928daa4dc3391d4731aebd7824b84fbb89230a52b3fad066727
size 54189
