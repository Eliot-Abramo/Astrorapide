version https://git-lfs.github.com/spec/v1
oid sha256:9691b8991c58a1907d9f846c4c8a48cfb76251aa3fc9f89f779ff0998030393f
size 13362
