version https://git-lfs.github.com/spec/v1
oid sha256:91a490b9166c8d2bc279124c1dc05dc9f9d48a58cb0a5b5fcb48b7577d479353
size 14531
