version https://git-lfs.github.com/spec/v1
oid sha256:e30bef57926186f2c06e6cf602d2cc84f92376a8b9f2be1f53e34a107f94579c
size 76095
