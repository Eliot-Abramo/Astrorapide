version https://git-lfs.github.com/spec/v1
oid sha256:79632b8c32378820ec0ee96530555989e4dce5397ac8017a47dc2b499c381887
size 7274
