version https://git-lfs.github.com/spec/v1
oid sha256:913e97eca8b56c2ee5b56576602f33b0d3568275a29592778020c894c0f2a3d9
size 54967
