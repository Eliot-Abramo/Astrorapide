version https://git-lfs.github.com/spec/v1
oid sha256:81db5439ddb51cafa5498ea5b35657044350d90905117adef22f0af3b93ed086
size 126213
