version https://git-lfs.github.com/spec/v1
oid sha256:e2a24e0ab6434a7389d5523f841585f6797328eeff39178052191a4afc3afc5b
size 2118
