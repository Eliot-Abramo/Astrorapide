version https://git-lfs.github.com/spec/v1
oid sha256:21ea951ae622a36f0498fdb9f325c25c092f9ead019e685f9768511e3aeddd82
size 2426
