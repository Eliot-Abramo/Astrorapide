version https://git-lfs.github.com/spec/v1
oid sha256:fceac50839a6f3c8f375423902a523e7fbe161a15753b42b21cdd7e8189d1ea6
size 1889
