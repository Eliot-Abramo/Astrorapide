version https://git-lfs.github.com/spec/v1
oid sha256:b349b5f0c2585766ea1519f1ba60b4ba8d58884d39c62a20073fd48a2a0590d0
size 4491
