version https://git-lfs.github.com/spec/v1
oid sha256:47aa1c08ff1fc4d980615cea34c2179c7e39e65ac09b9019e561c11dc7fc35ec
size 92653
