version https://git-lfs.github.com/spec/v1
oid sha256:f258c1bbc6c3c56c7f41e51c3bf288ffac67fe316ab6b6533e5782a10244821c
size 44495
