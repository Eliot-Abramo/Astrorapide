version https://git-lfs.github.com/spec/v1
oid sha256:f2b78ce8eb378c44f59830508bf8279751ac74f9ded6cec29356c9e96db58a2f
size 3093
