version https://git-lfs.github.com/spec/v1
oid sha256:9062b9ed7bdb85b19762dc057338a2079cc0ee6c4f6c37d45d1fcf837fcfd0cd
size 43398
