version https://git-lfs.github.com/spec/v1
oid sha256:fb26e8da1a9a4a5faf505528b3695f0ad91c72138a9c595edfdeb6e31940a6d0
size 24470
