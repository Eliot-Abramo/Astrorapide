version https://git-lfs.github.com/spec/v1
oid sha256:1fd3a73b9c001b6de0029e2102b547ead3c329baad256bd8610f0ccc3e0eb0d1
size 54961
