version https://git-lfs.github.com/spec/v1
oid sha256:c5881dfe6b394061eaa6f0a7c8b6f6ceefc658bfb0c1f4a5a5a2a82dd36dcefa
size 5542
