version https://git-lfs.github.com/spec/v1
oid sha256:a9fdb579acaa7587a509775204c96dadc51eb28382d50a5dc459cfd4727061ec
size 43952
