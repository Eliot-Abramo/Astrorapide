version https://git-lfs.github.com/spec/v1
oid sha256:d1c38791b69638a2faf4ff210cd04eb4ef496a323976a6c2e52f0b8edb68fd5b
size 54818
