version https://git-lfs.github.com/spec/v1
oid sha256:0e10476f1d61b58a8526247456b6557396106a1551b2a81ad0e7913ca8394cca
size 14527
