version https://git-lfs.github.com/spec/v1
oid sha256:227b02880cf19c72bacfed23b32c221acbdd0003c78ab5ffc2056f394c72d6ba
size 47885
