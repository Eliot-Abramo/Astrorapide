version https://git-lfs.github.com/spec/v1
oid sha256:b399b0eb0ac26b60f855c1c5d89afc4c8a6002aae0dfef0854446a26484a3aca
size 40268
