version https://git-lfs.github.com/spec/v1
oid sha256:ce12e3d0207717378182f01320d81ba2d748a90966055e659757ffe33e611ce6
size 43934
