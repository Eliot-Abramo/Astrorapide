version https://git-lfs.github.com/spec/v1
oid sha256:877fba90596611db19220058ca34b62dee58a9dfc06972b4a625e89292088ee1
size 2091
