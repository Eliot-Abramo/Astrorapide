version https://git-lfs.github.com/spec/v1
oid sha256:32ff96f731872a913796eeb655fc3fc17e03c6742f48f247ef49967a16c57f46
size 105228
