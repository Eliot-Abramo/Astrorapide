version https://git-lfs.github.com/spec/v1
oid sha256:34ae1a6362e1b382c28a18ca61d382b6532d7ec2f37f4600b69c1dbaa8a463f0
size 13387
