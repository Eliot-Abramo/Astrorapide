version https://git-lfs.github.com/spec/v1
oid sha256:d852f4c0df8c676f66ca26858b55737b26bb743621049691c4339ad6c22a943b
size 2108
