version https://git-lfs.github.com/spec/v1
oid sha256:dac61bdeca002715dc0d56d6ef5756d8d3638be5ea17bd2b2fda008b2558e0a0
size 41264
