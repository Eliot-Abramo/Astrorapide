version https://git-lfs.github.com/spec/v1
oid sha256:759247eb21eabb5962b546b24039d0dd1d1c4a32f17d6040bd5271a4eae27f1f
size 9287
