version https://git-lfs.github.com/spec/v1
oid sha256:5a0da1dbb13139d3440ccb350689f93472c800c515e0a4463445e49caf2b9043
size 54893
