version https://git-lfs.github.com/spec/v1
oid sha256:146543679375ad680f950eb37af48ad71e7299fe35156ad9c47906dcf200ab8b
size 17623
