version https://git-lfs.github.com/spec/v1
oid sha256:3e8290e84b07bbdf304df817219476b619df7f880101ce90454cd37f09306b87
size 58277
