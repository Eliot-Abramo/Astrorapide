version https://git-lfs.github.com/spec/v1
oid sha256:f669bc486417315653c4285bcc580ec087c922a941f6d927732b3a46d74a2ca4
size 14339
