version https://git-lfs.github.com/spec/v1
oid sha256:932655eec0dde46eaf47dddc039dcf8b1f5fc02814362c38b057e98269490837
size 13370
