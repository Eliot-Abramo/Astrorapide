version https://git-lfs.github.com/spec/v1
oid sha256:233f5ad7387120f6a91b10e11d1bb7bd247d0f730c156bc2b15026762380b675
size 10650
