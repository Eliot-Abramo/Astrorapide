version https://git-lfs.github.com/spec/v1
oid sha256:a244f4830e3969e1f5524487e1861cee11c99423ae9b8216dc2562b480f74bca
size 2054
