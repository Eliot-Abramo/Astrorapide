version https://git-lfs.github.com/spec/v1
oid sha256:2896c8109298b71b2e4bca44bbd57fb89a4ce33e75c9af3a463d114523976008
size 2825
