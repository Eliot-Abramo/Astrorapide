version https://git-lfs.github.com/spec/v1
oid sha256:d220107988c58163c578bddec6f6a4580b926fec96743c2c8737bede5bc43e76
size 3103
