version https://git-lfs.github.com/spec/v1
oid sha256:888e26bb15babfbe8cbf344a6745a26d0b07a3190507d5213d134cca82865a8a
size 26490
