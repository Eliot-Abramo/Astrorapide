version https://git-lfs.github.com/spec/v1
oid sha256:2f8e4b0480b852bcd7c42b35e9bfb89501a28e7f37bcfb725db941c0af8d3c72
size 2401
