version https://git-lfs.github.com/spec/v1
oid sha256:8a40c766f7e85af4994362079cb96ff73ec748afb61494322a97e5d74268ab97
size 10113
