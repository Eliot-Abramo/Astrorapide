version https://git-lfs.github.com/spec/v1
oid sha256:a8aa6f696d17c9cd61a91f2a24630043bb5ecb1bc539b26e509c921ddbec8583
size 2082
