version https://git-lfs.github.com/spec/v1
oid sha256:12ec7e38c6d8d7322e5a177992c1c553209133eb631faacd0102a1c33b38de3c
size 9225
