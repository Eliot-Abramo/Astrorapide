version https://git-lfs.github.com/spec/v1
oid sha256:72eae43abc0a58502869dfcf58f6bfe63737234c23e4cc19d6d6eda2339fd510
size 5257
