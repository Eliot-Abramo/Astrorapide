version https://git-lfs.github.com/spec/v1
oid sha256:36fe1a7a196cddc1e5fed483ca91cea7d941f03c614c1463e6ba72fc37e85ecc
size 3107
