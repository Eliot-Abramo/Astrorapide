version https://git-lfs.github.com/spec/v1
oid sha256:aff8910d47bb358bffa03d34f30a49d187d98cc28aca02abf95cdf1d9aa62dd6
size 2112
