version https://git-lfs.github.com/spec/v1
oid sha256:50444f215b0bdb693cf7b326adc887ed4d48e10458aad84a1dd139f71fe2414d
size 19855
