version https://git-lfs.github.com/spec/v1
oid sha256:894ddcb41f24f74b948c2170d320c7c85f59d5f2d7a1b04a091b4a681fd34dc2
size 5380
