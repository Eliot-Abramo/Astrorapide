version https://git-lfs.github.com/spec/v1
oid sha256:1d9d77832c5423fc066ea88e7e16543b714bfe4c727e57590fab5b2c9d45000b
size 2110
