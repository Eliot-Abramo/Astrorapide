version https://git-lfs.github.com/spec/v1
oid sha256:e3209d23864aa37abd892d43041e89b2a3ce742788579024376cd257cf054649
size 19829
