version https://git-lfs.github.com/spec/v1
oid sha256:73201dfdcb9eab49a5464914f2bfac6ac286ba358301d421dc7ef49180549d15
size 2092
