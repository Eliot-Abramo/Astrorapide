version https://git-lfs.github.com/spec/v1
oid sha256:13e7c682da0d58997eec486d8c243f99458f2a1271e5cb6b7ef5d65ceea4e5e6
size 54997
