version https://git-lfs.github.com/spec/v1
oid sha256:f5725e475b7db1ab9ff4072159305a45ddaf9ebb8bd996b8ba7e9b580ce77c1b
size 2839
