version https://git-lfs.github.com/spec/v1
oid sha256:5fb38f9e359fc8dc87f7aa8385b4f11a1e92a4f6d8058fab405adcfcbe7a0702
size 216928
