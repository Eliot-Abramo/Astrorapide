version https://git-lfs.github.com/spec/v1
oid sha256:01f0a67322bb2b628b8f116719d8f309ae42be0484ad0634b08bc29cb9514557
size 2839
