version https://git-lfs.github.com/spec/v1
oid sha256:133f0993425bacb02f6de8ed5e0ad3c1b648e059b3db6e5d47cfc3e4518bb3ea
size 5313
