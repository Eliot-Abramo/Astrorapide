version https://git-lfs.github.com/spec/v1
oid sha256:980d3e153c18d8042a64dc6acc887049c35848ae6509b9fbcb053a3dfdba745a
size 13401
