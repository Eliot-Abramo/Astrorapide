version https://git-lfs.github.com/spec/v1
oid sha256:6211af7b14e181513990f019078dca85e5d90a25900e01402b688ce79609026e
size 54817
