version https://git-lfs.github.com/spec/v1
oid sha256:d41e8aca0d48a111d87eb32c55c391e5424e6dcb033d1ac350e0974516ac6a4a
size 48847
