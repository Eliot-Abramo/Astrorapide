version https://git-lfs.github.com/spec/v1
oid sha256:0e8124f09577097b2b49b5a08d0cdf81b227bfaa6b828799a9989ecb9e3913d2
size 1837
