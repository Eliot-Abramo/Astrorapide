version https://git-lfs.github.com/spec/v1
oid sha256:dd525905ac33d9d66b8d8355b61bd41855eec6ae741d7eaa0a5d5d063939d47f
size 13390
