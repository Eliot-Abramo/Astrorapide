version https://git-lfs.github.com/spec/v1
oid sha256:120c570049dec4d6aea0a7d12766311451aa6d088edc278ae9b28a738ec0562e
size 5313
