version https://git-lfs.github.com/spec/v1
oid sha256:c83735707e4ddf9b85d8ab18932971c335ecdf8b3d6156d8a551acd1b9974c3c
size 17613
