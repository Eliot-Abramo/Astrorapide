version https://git-lfs.github.com/spec/v1
oid sha256:a239f8aa9289c09f92ce4c8e7e96ec1cd2c8e4a9fc83c2c06827af2964a9ba39
size 43952
