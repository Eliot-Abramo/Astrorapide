version https://git-lfs.github.com/spec/v1
oid sha256:7ab6b41d0c676e76584c45804b6ee8eefed8d079443552061b6ef00506086dae
size 4477
