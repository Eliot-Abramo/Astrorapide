version https://git-lfs.github.com/spec/v1
oid sha256:87431b29a7cac86a0e0a18fb437aeb7b61d1f8ca0e6ff38f9d160f23c0804dd1
size 17900
