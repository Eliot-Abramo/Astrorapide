version https://git-lfs.github.com/spec/v1
oid sha256:e07a30932bc755f6277b158355cfc6266f25dd857ccf99ed7391aa41df87b397
size 83239
