version https://git-lfs.github.com/spec/v1
oid sha256:3f9d77e1857e803131f54254fa02ef295d3f35c35ccf2beec9ec7a44994c1f67
size 2104
