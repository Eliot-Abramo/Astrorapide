version https://git-lfs.github.com/spec/v1
oid sha256:38741d241438a39940f81448225ba2258009fb3db072f076f7a765819dec902c
size 5313
