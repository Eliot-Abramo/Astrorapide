version https://git-lfs.github.com/spec/v1
oid sha256:658d7df405c356ae5558d59541742145d5e2db51b1d9809ffb2a4864b08cb374
size 17638
