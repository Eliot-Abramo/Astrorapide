version https://git-lfs.github.com/spec/v1
oid sha256:0df098cd9e8bb430d5d872ba3ce181a26af1acb3652d4596da5dd0fed7aaea62
size 72470
