version https://git-lfs.github.com/spec/v1
oid sha256:8b5c0addd381cd9d8599af872ba3849c5f9616bb91e1af3b5d8dc7adead03f7e
size 2112
