version https://git-lfs.github.com/spec/v1
oid sha256:371015f751908ad2f523fe059c8efc2332706fa675ce51448a5e37c4d3383121
size 13034
