version https://git-lfs.github.com/spec/v1
oid sha256:3f63fb977607e4f40003673b468d4e53a3566895ef57ccb02ec8745527265476
size 48772
