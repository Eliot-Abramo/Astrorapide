version https://git-lfs.github.com/spec/v1
oid sha256:f4e889a0dc3f2126aa47b3c17f043b467bd620546212d64b1ccdd17c185d2514
size 76095
