version https://git-lfs.github.com/spec/v1
oid sha256:4a85db92bc57dd0820dc8f05d479ec5272d7efdb5d387c78600220c25bb2490c
size 129616
