version https://git-lfs.github.com/spec/v1
oid sha256:5935d7c889da66e787d23269bc08223df3d0f4528b6ad76fecc8c0ba98bde982
size 5531
