version https://git-lfs.github.com/spec/v1
oid sha256:3af69e8dd75694115d0c99924a27eed152b18e38e68128485ef15d2c5856e05d
size 2112
