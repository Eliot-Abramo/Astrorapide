version https://git-lfs.github.com/spec/v1
oid sha256:c13f377e68ad628ecb0551ac00257cadc84334ec290650742a69b4a66ea365e8
size 14524
