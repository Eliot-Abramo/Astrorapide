version https://git-lfs.github.com/spec/v1
oid sha256:a0366ce5b7691a05282e5fbbc5629007918b4e5d7abd16ca697d3a3398bace11
size 12940
