version https://git-lfs.github.com/spec/v1
oid sha256:c8915928b751c1251afd602a56be61335ddb0859d85453699c862bdc1a2f7b2c
size 5486
