version https://git-lfs.github.com/spec/v1
oid sha256:25b58faa04224fdb846f6ee7eca1454226faa2a93aff15f6f4d79b0f54e6a159
size 20978
