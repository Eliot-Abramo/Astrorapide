version https://git-lfs.github.com/spec/v1
oid sha256:ee3bb9481fb15a3c6ab82cf968b33b4eae4747858486e5445144e2e24848ded7
size 46282
