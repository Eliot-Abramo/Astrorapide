version https://git-lfs.github.com/spec/v1
oid sha256:95549cfa98c164fbe4ceebd03e75365141ad8734c5cb58ba2d6caae2afd08eae
size 3093
