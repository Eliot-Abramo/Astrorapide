version https://git-lfs.github.com/spec/v1
oid sha256:1a0fb05fefc6047c92d3810663c2c5995a53e72d1716e5bad98164cff5daa0b0
size 2287
