version https://git-lfs.github.com/spec/v1
oid sha256:4e69a22928c61c05da4a56b59f8dca66918db3e841cc7950fe3edc33969c7aa4
size 2092
