version https://git-lfs.github.com/spec/v1
oid sha256:f6d129584023d2ba9943f10ab5f29b5c93b3c26b4845041b1ba86ac117f2c210
size 14658
