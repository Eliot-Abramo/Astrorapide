version https://git-lfs.github.com/spec/v1
oid sha256:12eace44f6d78452528ddd6b21d1772c31a8ab52398d4b8cb27d1cc384670a43
size 17398
