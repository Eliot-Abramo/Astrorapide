version https://git-lfs.github.com/spec/v1
oid sha256:16d5130dc97c1e8dac545532f102a89bd1acc963f5e958295e6fd9fa04824e22
size 113822
