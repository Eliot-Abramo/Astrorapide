version https://git-lfs.github.com/spec/v1
oid sha256:4ef1d3a7b5140c548bb7a3218ddadc07a5595c2bffcede6ee7ca8779dd824b72
size 13177
