version https://git-lfs.github.com/spec/v1
oid sha256:3035a8afa06d73bd65f586e00bde10b331b60af3a83d1435b756d0faf3d53677
size 54873
