version https://git-lfs.github.com/spec/v1
oid sha256:757ffa01bc54f8397d0db69c2d71bf8a032b945ad9e14b2b67cd7fc8acc342a0
size 76095
