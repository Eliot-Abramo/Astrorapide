version https://git-lfs.github.com/spec/v1
oid sha256:50fc59c04a2a3a94c3dac97a29e0d64490dc5efbd10f075f2a59dd0146e6271c
size 2118
