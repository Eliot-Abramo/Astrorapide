version https://git-lfs.github.com/spec/v1
oid sha256:488e9224b4293d8f7d223423cad0e1d8b3f7ffb86c2ccb73a6d829e2d8804d12
size 14532
