version https://git-lfs.github.com/spec/v1
oid sha256:232cc7991c85c2d434b8003436b191636f70977f2fd6fe059282b31c72f67ff4
size 24472
