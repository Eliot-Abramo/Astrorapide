version https://git-lfs.github.com/spec/v1
oid sha256:852a3c6ebf132b6c95940aec182492801013e4e0e002c213bcc964aa8f18fbaf
size 12510
