version https://git-lfs.github.com/spec/v1
oid sha256:871df307d33d103ef6e1d1ea18e78533ae4092849cbeb8588522216b40f5372d
size 39729
