version https://git-lfs.github.com/spec/v1
oid sha256:714cd01710bc407effd72f80b288f4741398fc6cfb59a7cb34a3709defe41dca
size 1508
