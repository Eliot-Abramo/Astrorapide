version https://git-lfs.github.com/spec/v1
oid sha256:584853ece815741e07e8f116b7879ec856812d2ff199239256e501a38e3f8c5b
size 46402
