version https://git-lfs.github.com/spec/v1
oid sha256:488f6512c7782bb9c4fb80074502027f75709d2d9ee26997e1306b573eeab32a
size 14532
