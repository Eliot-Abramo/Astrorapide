version https://git-lfs.github.com/spec/v1
oid sha256:cbebcd30c1aa046677bda5a208acd2412e61e7ee831f1b81b7baabb9f843f17c
size 2426
