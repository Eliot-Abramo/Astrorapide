version https://git-lfs.github.com/spec/v1
oid sha256:42ca6cc847e5e5af9b27dab9dab99432366f2c1aea0cdab6eb4651a9441fb85b
size 4254
