version https://git-lfs.github.com/spec/v1
oid sha256:2030cbc4d6662bea492edba3d45a9a201a6123226498fea677932e17f9f6b1e1
size 76127
