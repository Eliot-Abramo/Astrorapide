version https://git-lfs.github.com/spec/v1
oid sha256:eeb47126a7a3f53f29d839426a666ebb7749aa420d76947f582a534c23bf8d71
size 24272
