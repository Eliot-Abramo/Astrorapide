version https://git-lfs.github.com/spec/v1
oid sha256:b406522be2206628dc9fe05734871a0110401f4a7bd4bbb04c0f691497f43794
size 19571
