version https://git-lfs.github.com/spec/v1
oid sha256:9c3f3c99e71116fd7a715b14bc74b09ac994c0b36a332796554398f31a55ea2f
size 3979
