version https://git-lfs.github.com/spec/v1
oid sha256:d3502b1480909c6e14ab375b38c186cbfa0e97cebf9ae14ff1284f9f378b1d99
size 1903
