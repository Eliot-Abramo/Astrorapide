version https://git-lfs.github.com/spec/v1
oid sha256:e48475ecb2b02b2fb25c0fa2b3665fb612c9b92762f82d1178afb8a9ac000085
size 48202
