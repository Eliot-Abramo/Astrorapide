version https://git-lfs.github.com/spec/v1
oid sha256:d66c16fdf2c9be28085a99063b7d077d94902f84ace29d4307e1642b7fc7ca3c
size 39060
