version https://git-lfs.github.com/spec/v1
oid sha256:03b80d7973cef94380321af054e2ab393907a47bbab0d14dc599c49168b40fab
size 2094
