version https://git-lfs.github.com/spec/v1
oid sha256:222c1b35a2cf113560df35bb75a5152c798e93935bfb87d6740d4aa94b48e836
size 2004
