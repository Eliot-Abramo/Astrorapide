version https://git-lfs.github.com/spec/v1
oid sha256:067fc6b421eb4f3dc08fe27e3750b9665bfc1228561325b8d5072f5ca263807e
size 2413
