version https://git-lfs.github.com/spec/v1
oid sha256:29cc2eb8f4b4c0e68fb4757ad6d331a139650d1e22c92f0fafb837d4cd66f26d
size 13459
