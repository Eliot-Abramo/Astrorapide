version https://git-lfs.github.com/spec/v1
oid sha256:c91570be5ee6a91c46279eec4babf42e222c3a58cc7174484471cb88ddfb51a7
size 17651
