version https://git-lfs.github.com/spec/v1
oid sha256:45c6f8f8c0b6e02a6f875398f52fb87d01fd30dbaf93245967ad598ac029fcb6
size 92389
