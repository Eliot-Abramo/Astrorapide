version https://git-lfs.github.com/spec/v1
oid sha256:e08c2a7147724ebc0842aaf6e8c487bf3a3d21976bdb9ef9655674f6f4153921
size 13235
