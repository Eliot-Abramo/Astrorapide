version https://git-lfs.github.com/spec/v1
oid sha256:9ab6de85de123a1f3e26ef624dbec4a2f7c81dbf8116b78170deb7a0968c391f
size 10099
