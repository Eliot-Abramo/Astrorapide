version https://git-lfs.github.com/spec/v1
oid sha256:8fcb24053ddbcb86be4bc4a49e6e94aa25b02ae0328cdf2c984d33ba20f70c15
size 12506
