version https://git-lfs.github.com/spec/v1
oid sha256:a622ccaf5b1c4a97996aba6526d7ff601cbef06460016850388c355dddc19d68
size 13376
