version https://git-lfs.github.com/spec/v1
oid sha256:953330d1c2158b75275ed7bcb82ee3e6cc6bb40d1eec70523dc4bb3fde7b558e
size 6234
