version https://git-lfs.github.com/spec/v1
oid sha256:2eb89e47d3b5463ee42161692ad111c31abe11534d61fb0251f623f2d2e353b8
size 105228
