version https://git-lfs.github.com/spec/v1
oid sha256:a420c3f62cb48d0b321407d92ab909c6ca8bb0a91761ce632e0a757b8fe6ac26
size 13414
