version https://git-lfs.github.com/spec/v1
oid sha256:43b5caab9b55a5355a8fed0a4b82d86439616bdf2f3ebefe22fd2ece1abb7c36
size 5321
