version https://git-lfs.github.com/spec/v1
oid sha256:89b560111c2e5489944c7298264d9fe42fde787f1698b90fbc4f8329064777f6
size 2840
