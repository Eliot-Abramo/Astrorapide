version https://git-lfs.github.com/spec/v1
oid sha256:388be5beb34d9ecdedcc88d3770b993cd8200fb42e0a3ac22f3d2c2d83231e8e
size 38448
