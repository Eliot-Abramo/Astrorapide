version https://git-lfs.github.com/spec/v1
oid sha256:840935a185266ce553715b0962fbed5d980afe745efd33e9c8931a17a3103b07
size 146473
