version https://git-lfs.github.com/spec/v1
oid sha256:3813bd478c57c0274b392a8a6e968a7289bbaa675702b084cdb5a02f759a45d6
size 39679
