version https://git-lfs.github.com/spec/v1
oid sha256:b0b12f65482b6b77d2af4f3ddd63c20fdf1a2ff220ddef4614262fb4307038f2
size 39166
