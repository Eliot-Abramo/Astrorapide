version https://git-lfs.github.com/spec/v1
oid sha256:9d9a92cd692c311f46fa2e3cdaac759d7269c93913483f116037f2c118e3ef08
size 17692
