version https://git-lfs.github.com/spec/v1
oid sha256:b73ba0fd83cca07486c4a482698873bef2a0415fb6d14b27261a04b513b249cb
size 20978
