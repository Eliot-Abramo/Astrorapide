version https://git-lfs.github.com/spec/v1
oid sha256:1099107891cee64df1fb55df87f186ff1ab29e8033980b11caf9464bba22e54b
size 24472
