version https://git-lfs.github.com/spec/v1
oid sha256:678adf45a243714728482d2d0ce8ed864eef66ba3198c9b712bf97ad3a8382b5
size 2837
