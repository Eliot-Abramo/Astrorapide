version https://git-lfs.github.com/spec/v1
oid sha256:a4cb21aaf9b04037460d782f62e7bb257c73fab286b8b824442571ac8120f888
size 106755
