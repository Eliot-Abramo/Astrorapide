version https://git-lfs.github.com/spec/v1
oid sha256:5be7a0ea7e82d9cc78fd4ef3fde71fac3b85c2bc8a8816b8f76f6e8933091c2f
size 5313
