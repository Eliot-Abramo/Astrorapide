version https://git-lfs.github.com/spec/v1
oid sha256:1446748e6b01e1fb4924ddd7d23cf229a8dd0a2adbd090b354bc9bf8aeb8a46f
size 38503
