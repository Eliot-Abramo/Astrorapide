version https://git-lfs.github.com/spec/v1
oid sha256:a57d5e9c3c4a56cddb62f796e0ab2dfa1f3c2ba039c6e9a1578fe802b4516ff1
size 25758
