version https://git-lfs.github.com/spec/v1
oid sha256:747eb763c154f5893f8441a133651a4438d10517f81c8bf193428cd14e2c512b
size 2086
