version https://git-lfs.github.com/spec/v1
oid sha256:41805bd3084c12dec1949d6a01e60bfcdfef2d547cfb1f59e8ee6fc4ecaaae1e
size 24470
