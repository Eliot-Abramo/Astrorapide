version https://git-lfs.github.com/spec/v1
oid sha256:7c2de7ae847ef624869dcb6e0cef7ebf2c824945d255ab52754854370b998f32
size 2401
