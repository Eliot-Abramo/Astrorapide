version https://git-lfs.github.com/spec/v1
oid sha256:186bb6c2464c19668d32b3da779252f61011105259805d5e40c6cd14a42dd72e
size 6264
