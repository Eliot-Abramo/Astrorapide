version https://git-lfs.github.com/spec/v1
oid sha256:995a50bbbbab92525d090ca824cca2903b67dbe3ba7095ca13f88683283a0a42
size 53713
