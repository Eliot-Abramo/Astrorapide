version https://git-lfs.github.com/spec/v1
oid sha256:04770b61e36be8416a1a54e1d2103ee73d9754a570f672bb70496ad5b68c5b89
size 1903
