version https://git-lfs.github.com/spec/v1
oid sha256:a56fc87312598ec1b5d08596c745676304cee3c885c192c1989d3e7bdcfecefb
size 76095
