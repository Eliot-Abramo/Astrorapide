version https://git-lfs.github.com/spec/v1
oid sha256:e4a49b841aa75f5f5ebf8758d317257cddf66b78f7cf3685a77de2d0495e186f
size 20987
