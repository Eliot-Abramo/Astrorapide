version https://git-lfs.github.com/spec/v1
oid sha256:e8907289167cdfe7643e9ed136dbebaa0a236338d76adb56e4a70181213571b3
size 14658
