version https://git-lfs.github.com/spec/v1
oid sha256:c823127226a7ba75bf227950667bbf5ca857ca8a1766cd32becee42cd140b489
size 2110
