version https://git-lfs.github.com/spec/v1
oid sha256:6ec9c3c424390835206d60160a8d10f4dd2eb3d318a6b440e68158cee5d603c4
size 82870
