version https://git-lfs.github.com/spec/v1
oid sha256:e5b41da0675f9e5899dc032a9300da1ef32c90a5f23264bbfbce9f6a1c7e9ce1
size 18135
