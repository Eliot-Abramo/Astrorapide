version https://git-lfs.github.com/spec/v1
oid sha256:147d980c5cb8363cee7145f342dfbfb3d6e669d924a3b42a7324590c0e81eb30
size 20987
