version https://git-lfs.github.com/spec/v1
oid sha256:c90624533dbc2ff671de2d54c80b1d4e095edd09ba4657b461a864f25f751bed
size 17947
