version https://git-lfs.github.com/spec/v1
oid sha256:04eb58dfa1ee32f2045d334043222d683a4a6889ae9f4e73923d29529280b745
size 2415
