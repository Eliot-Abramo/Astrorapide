version https://git-lfs.github.com/spec/v1
oid sha256:1738b13832aa9c8a5ddd53d74a23f9168b3d99965c2dc5c354eaf9f67e2c27a0
size 13407
