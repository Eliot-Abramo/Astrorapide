version https://git-lfs.github.com/spec/v1
oid sha256:764f55f86998c8296bc65d664a63c8e250ad1ed588c3f455166229914f6b5cc1
size 40088
