version https://git-lfs.github.com/spec/v1
oid sha256:cccba014ad900e1b6e248aafe1cd5180b1e7f5db7f201b6dca34e8817ebb298b
size 61359
