version https://git-lfs.github.com/spec/v1
oid sha256:57c73d251b6f1759a79dcc3de3d1feadad39d0a8a66e099155ce16b7e0aec0b4
size 2106
