version https://git-lfs.github.com/spec/v1
oid sha256:ad085e16965c4dcfa8200723386b612638f2abc9c0e75427849045fc759ab405
size 2093
