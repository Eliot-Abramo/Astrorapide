version https://git-lfs.github.com/spec/v1
oid sha256:4bedac9e020ada0d098b62e295ab4ab480caccb688b275de8fe87149aceaa927
size 20970
