version https://git-lfs.github.com/spec/v1
oid sha256:9576b78088a58941c75541d8aca7b2c129aaa28aaf94471fca9178830b65319a
size 56368
