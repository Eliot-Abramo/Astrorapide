version https://git-lfs.github.com/spec/v1
oid sha256:c69d6d891a47aa0f60ed7dc890f7c818ee337d8cec18d7c42e3e22b0913940ed
size 2118
