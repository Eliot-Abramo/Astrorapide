version https://git-lfs.github.com/spec/v1
oid sha256:4813faa6d7b2b0a98a5dce12083c2d94853f7061536d3e707b5fa560a50298df
size 36092
