version https://git-lfs.github.com/spec/v1
oid sha256:9b2f1b87af155646dcb7a698170df81fe5654b316b3fcd2708b53158846da927
size 1899
