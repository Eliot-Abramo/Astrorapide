version https://git-lfs.github.com/spec/v1
oid sha256:4336fc401a80222b66f3ba1f4e744ecc321ab39c91828f6ac6f2e7389445c33a
size 43400
