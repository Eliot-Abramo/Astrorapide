version https://git-lfs.github.com/spec/v1
oid sha256:1cb2a96062eda31518ab20d760925d356bf181f4329c41f28479b36d37b98368
size 15713
