version https://git-lfs.github.com/spec/v1
oid sha256:ee746d02281a10b7ab48298b609b4c95588d061b127f3f2962beab9cd5bc49d3
size 13169
