version https://git-lfs.github.com/spec/v1
oid sha256:0ff9aeb979edc0c31be63b8e7ec4c14ae7e055ef1073d9d3e7212e3179b13374
size 105527
