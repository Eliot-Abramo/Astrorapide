version https://git-lfs.github.com/spec/v1
oid sha256:185e30e461a69443d1452deaeeb8810f8ee0d3b754207fe336d604c05c7e347e
size 47140
