version https://git-lfs.github.com/spec/v1
oid sha256:25225a0dae5bca19ec19a3c22262fa30552e075c9f0df57a5995cc963fb13110
size 10110
