version https://git-lfs.github.com/spec/v1
oid sha256:437d6e9ea61c5306a6a5367451deeb8e5015905ea150a94a365f6f39ad96fd78
size 39757
