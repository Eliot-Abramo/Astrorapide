version https://git-lfs.github.com/spec/v1
oid sha256:a6368d7b8f9a38c13ea46f56be42e596030162f000618ff0a36d163c0a84372f
size 2840
