version https://git-lfs.github.com/spec/v1
oid sha256:8b0c841ccaa6de480123c486e90aae5eda441aa550e348e728752eecbbfd5efe
size 47019
