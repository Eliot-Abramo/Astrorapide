version https://git-lfs.github.com/spec/v1
oid sha256:c13567e509748766d424afda9a3df8401ee298df9e4c68c726790dbffaa1c75f
size 13180
