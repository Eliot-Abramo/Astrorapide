version https://git-lfs.github.com/spec/v1
oid sha256:fec74f5febfdbe1d5fee8416cdea85d125268c76986ac6c4423459bb459284f3
size 9550
