version https://git-lfs.github.com/spec/v1
oid sha256:5a2e17c56a611ae09cf5fa495e89db41952fa35bc5b58eeb518dbd580bd90f4c
size 2005
