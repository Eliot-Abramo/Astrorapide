version https://git-lfs.github.com/spec/v1
oid sha256:1a550709d6db030115a9e64b539e8a8836ec09e85f67bfcc664b6c4514560fca
size 10650
