version https://git-lfs.github.com/spec/v1
oid sha256:0a283312121047ec079b86a14f57168016ae435c90aa257a391bd87a447b1469
size 4489
