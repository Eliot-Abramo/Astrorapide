version https://git-lfs.github.com/spec/v1
oid sha256:01d93b58af1d7add115f9b7177525cfcbda3719e227a1c14811a735e77e75b91
size 3937
