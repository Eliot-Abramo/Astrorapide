version https://git-lfs.github.com/spec/v1
oid sha256:d45158ed0ae33c912a7552cadb904516cf41213d42f5d455f1ad1d97f01cc5e3
size 34453
