version https://git-lfs.github.com/spec/v1
oid sha256:acf3b6487f01948eee87ad58e884e00ba08f92860af820efb3e78768373aaa84
size 13390
