version https://git-lfs.github.com/spec/v1
oid sha256:1431f1407cc11da41976c5b24d1aacf6ef5c5bb06e16bb2e17331f1383eb987c
size 54997
