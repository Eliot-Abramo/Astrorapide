version https://git-lfs.github.com/spec/v1
oid sha256:714476698acecb9b55069eaf9c0627a13fd64d549f94a0bb56c5ef0d5d5ca7f5
size 52690
