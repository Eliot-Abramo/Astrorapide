version https://git-lfs.github.com/spec/v1
oid sha256:5cb17b7fdf6a7415db3c708610fd9f2e9bbf3318b1e84ac7e6f96bb84d831481
size 12954
