version https://git-lfs.github.com/spec/v1
oid sha256:7ef333d2ff4fbe79eba61278ab96b756043cfcefe4cd3659c8b95ad84d01b171
size 43400
