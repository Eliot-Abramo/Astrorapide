version https://git-lfs.github.com/spec/v1
oid sha256:a24c6ad35705fd34bebc79ae184745b6ed57d0d98a0cb634f652c7f7c0476b18
size 13473
