version https://git-lfs.github.com/spec/v1
oid sha256:b0fff9d1308342eb808f333c3571e15a662841d4a846b9166b00f2efe89176f6
size 66468
