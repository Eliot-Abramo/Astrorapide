version https://git-lfs.github.com/spec/v1
oid sha256:51d05220957d626f951e78c81279e5833c58accc38f39bd529b22581ccc728f1
size 2833
