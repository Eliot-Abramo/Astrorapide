version https://git-lfs.github.com/spec/v1
oid sha256:28b81ab2dc56a890c6cade969cf6a42e8407c885051b7aee9e82959007f91a9b
size 66121
