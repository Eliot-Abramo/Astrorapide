version https://git-lfs.github.com/spec/v1
oid sha256:9782e8ffbdb8ce6fc70888b61b036aae9c33ae7906566c0cedf0c35771093cc6
size 2116
