version https://git-lfs.github.com/spec/v1
oid sha256:a7ffded1c7229a1381c7d3476c61e63e85bacf950bc9a4943db8a09a3e58776a
size 54179
