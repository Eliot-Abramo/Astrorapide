version https://git-lfs.github.com/spec/v1
oid sha256:f277f8dfa9ad103068c2f0e3cd6cda3f0e9f2b74c96c61b9d5d9509c3df9e105
size 2110
