version https://git-lfs.github.com/spec/v1
oid sha256:9790ef64f601e5ff38bcf09c7e376b989123e46c2804628b686c497f76487ac7
size 14656
