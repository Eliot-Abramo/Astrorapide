version https://git-lfs.github.com/spec/v1
oid sha256:f407e3b7955e71a6b44322936ad110ef8aeb39ab8b79f06bc92e6e14b2a8f334
size 10147
