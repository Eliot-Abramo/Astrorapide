version https://git-lfs.github.com/spec/v1
oid sha256:495c7420672fd31ef1a54e7b21a338ead2f0830541e4a3369c5210f2dbf2c861
size 2426
