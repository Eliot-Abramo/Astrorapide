version https://git-lfs.github.com/spec/v1
oid sha256:b6ad5e826d7e9a54eb94a430972389cd87c22723301ba5f460e776893131142c
size 51592
