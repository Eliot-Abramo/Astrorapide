version https://git-lfs.github.com/spec/v1
oid sha256:963dbfa6bb9b5daa24e161668432a9a218c41af4a5858a4cc2b803992a70abd1
size 47899
