version https://git-lfs.github.com/spec/v1
oid sha256:7447a2a520b0cfe6935980c42ee3e7cc87f60a43fe0d4080b976d060cfd74b3d
size 5313
