version https://git-lfs.github.com/spec/v1
oid sha256:6493fdc077a1add62c1e7ba8a8385cb2135f79500df9db1f4c4e0b08b5fd0403
size 492805
