version https://git-lfs.github.com/spec/v1
oid sha256:13c80058fbd3919430ad37f9e70a465b55eb5b970e09b5db541956e09b6b3f1e
size 14535
