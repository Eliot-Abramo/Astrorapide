version https://git-lfs.github.com/spec/v1
oid sha256:9b252aaad891c17862ace5d9fdc7c666a94dc00154cc4246a2583bbd997e4070
size 7274
