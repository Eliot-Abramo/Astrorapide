version https://git-lfs.github.com/spec/v1
oid sha256:f9e5f9ca807b588f572cd92bd78d0d34c1a26e8ec3e7e2ce0b8364a50e48624b
size 7288
