version https://git-lfs.github.com/spec/v1
oid sha256:9563454ae2f4a41c9b787799e1144f0443af75481f8454f61f18f4ef7f1f8b50
size 13393
