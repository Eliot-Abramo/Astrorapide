version https://git-lfs.github.com/spec/v1
oid sha256:b6999a4bf3aa746aca3edcc52863d451ae5187dd9b156b045c89b4d91c90fc1c
size 5265
