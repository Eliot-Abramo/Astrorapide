version https://git-lfs.github.com/spec/v1
oid sha256:28004ec40bb3f06ea7ccd26c16d879d8e93c91b2ab4606bef7bf5f7c83e712ed
size 40111
