version https://git-lfs.github.com/spec/v1
oid sha256:97bd0ffc27f4de6d73257a55f9b01de21c43547788e2d22dc2e50672df7b17bb
size 7246
