version https://git-lfs.github.com/spec/v1
oid sha256:0dae4908bba3047c4b0badf1a71f31542153fa5090a97e452da825052a414e90
size 2124
