version https://git-lfs.github.com/spec/v1
oid sha256:295670ef4fe60b41c82168ca421a7bd455307e8c10f9ee77b7aa70d89867333a
size 2411
