version https://git-lfs.github.com/spec/v1
oid sha256:ab8af0d557de39693ac66c40bf1ba38ae2e73606fbb00019fec8ad82b12a5912
size 2114
