version https://git-lfs.github.com/spec/v1
oid sha256:57999f4e8bcbe3892c03e802b30fafd472d554caa85b112fa589d12523d1d8d8
size 14494
