version https://git-lfs.github.com/spec/v1
oid sha256:0872b6739a7873f045b8851c07afc3e996cb17092d702fdc3c11ee376789f887
size 147068
