version https://git-lfs.github.com/spec/v1
oid sha256:791dfb13e13f45d38efe7c1d63e46a7d0ed928de121b3d42f89754579bdcbc76
size 17651
