version https://git-lfs.github.com/spec/v1
oid sha256:b3abc12e4ded034e375deba76bb6977217f26fdab6897b350a68a59d0d2addc9
size 2104
