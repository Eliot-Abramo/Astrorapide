version https://git-lfs.github.com/spec/v1
oid sha256:44a4849e539447fa3aa976ed3b32fe2af49db2c7b3881cc6fdf789093192500c
size 44497
