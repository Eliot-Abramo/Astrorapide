version https://git-lfs.github.com/spec/v1
oid sha256:c931a46fa5687836a73246a1c1da1677bc67e6c8378a52619bb9966600fa11cd
size 24286
