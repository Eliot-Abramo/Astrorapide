version https://git-lfs.github.com/spec/v1
oid sha256:216733378382267dd5b6cec6a488edaeb66185e33df9f7cb626c8c7552c0f0fa
size 2108
