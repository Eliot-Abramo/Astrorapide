version https://git-lfs.github.com/spec/v1
oid sha256:fe0c924eb0a6b983b540e6f092a482ef95d05a2ca2c0061a2ed1f201ed926499
size 36884
