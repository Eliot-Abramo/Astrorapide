version https://git-lfs.github.com/spec/v1
oid sha256:5403f1739046189e823be91d966430042dfeeaa5a96bb54bda5bbd6826557ac1
size 18533
