version https://git-lfs.github.com/spec/v1
oid sha256:e9fdf46ceff447e2f31fe2155a2e27b3a399f7785cd418ba089daac9a8f3f9dc
size 19855
