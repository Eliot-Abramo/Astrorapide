version https://git-lfs.github.com/spec/v1
oid sha256:7c04f31a92420c781672ee3375dacec83ad7b21f0cc726e504999187ced03dcc
size 2111
