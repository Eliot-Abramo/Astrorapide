version https://git-lfs.github.com/spec/v1
oid sha256:fc97c3532da762fd5f41e8b6e1479037fc1ab0e44cf5bb8f1e1be874fcc4ec27
size 113822
