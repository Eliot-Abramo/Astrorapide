version https://git-lfs.github.com/spec/v1
oid sha256:8e45fe4af7d574cd99c37632ac6e7ee670608daecd784f3ed90832f59ca96a21
size 14527
