version https://git-lfs.github.com/spec/v1
oid sha256:707b45d048828f6d2bdca4b304f2b1f1d2871fd970b4cb6e40a079868bf95388
size 50928
