version https://git-lfs.github.com/spec/v1
oid sha256:8f0b698a0ed2055bea89b598115467d3f4052e3b020ed0db867b255e4d75f96f
size 14531
