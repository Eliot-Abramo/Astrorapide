version https://git-lfs.github.com/spec/v1
oid sha256:6db9f698a3c7a73afa2b6ea31483840961f4d17a8ee65d8e3a1464942d37fd9b
size 2112
