version https://git-lfs.github.com/spec/v1
oid sha256:da301ce24f05a210f41424543aa3452ad929ed70dbb6c481a7fd180891f587e7
size 5948
