version https://git-lfs.github.com/spec/v1
oid sha256:2add484300a777efe7f389b02041dfa60760d00cc66002cedcb531d6b39c577d
size 14497
