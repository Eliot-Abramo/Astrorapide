version https://git-lfs.github.com/spec/v1
oid sha256:6b76a2afe81f26aa6e14aebc72b5236bfb8d9b4e1f1c743bf563479dab474f5f
size 5257
