version https://git-lfs.github.com/spec/v1
oid sha256:9432de9c163697f202083dcec361f5b68ca406947187a0ab0d9f2fdbd549eb5b
size 17664
