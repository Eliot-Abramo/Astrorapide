version https://git-lfs.github.com/spec/v1
oid sha256:2d999435f15f78552a0fb14f35f3f75afb008f0dedf1810d5f93bf0febfd03ac
size 11602
