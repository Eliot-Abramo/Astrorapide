version https://git-lfs.github.com/spec/v1
oid sha256:27db909411d705b3f0ef1b210d7fde588d9b97ec3d144317e305865059c55d34
size 83269
