version https://git-lfs.github.com/spec/v1
oid sha256:7c964cca22ae354f6bc540d740a1f85f2322bbced2f425b5afcfc353ad6b317e
size 20190
