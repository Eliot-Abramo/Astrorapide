version https://git-lfs.github.com/spec/v1
oid sha256:e1113f4d0f7fee6351d78a5c9a4f8a9673a22c52f6c7d8267cf6c1941dcfe918
size 10116
