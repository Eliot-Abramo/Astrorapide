version https://git-lfs.github.com/spec/v1
oid sha256:b9cfa03f02fcc9ebb9f1a22b8af25a6ca849ef9229d2366987138b22de7d6b86
size 19671
