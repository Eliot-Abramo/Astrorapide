version https://git-lfs.github.com/spec/v1
oid sha256:ec1b3903d51c423379338779b718b126e6c45666fff4198c3ff7001ab40b3b3f
size 12948
