version https://git-lfs.github.com/spec/v1
oid sha256:f9659add07978c6ea8f889b33cbc5a82e66c029ecf8b61193f3d79da83b4b061
size 16524
