version https://git-lfs.github.com/spec/v1
oid sha256:dbfb84ac709de98d9d57dc6840050e932a1aeeaac2e3c94cbce11188960ca1c9
size 76127
