version https://git-lfs.github.com/spec/v1
oid sha256:eef362bd7052f9efa09b54bfca6428812835a17bb7273e8b2177a9e678585f60
size 2106
