version https://git-lfs.github.com/spec/v1
oid sha256:6397ffd4481f9a654c1a56124ba842f812651c0ea03807743d3b1741b8f86ce0
size 9287
