version https://git-lfs.github.com/spec/v1
oid sha256:0158a96e69c054128e03a457d0173c48c1ed09e50c51bf200c484ea2359fe38f
size 54060
