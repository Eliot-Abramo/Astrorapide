version https://git-lfs.github.com/spec/v1
oid sha256:34ff68ff84d9b8349589a7f4c5ee0296b893233a849ae01be1ae1c23c3d34853
size 13398
