version https://git-lfs.github.com/spec/v1
oid sha256:8b017bad1e025fdb5b0e3297cd6f99142c08cc2f40ac401c0d54e9d43f8b767d
size 54540
