version https://git-lfs.github.com/spec/v1
oid sha256:894882e89651ace0f9241ca9de31c46b58d8e292d7f0b63c2a8eb20f8564f40d
size 14503
