version https://git-lfs.github.com/spec/v1
oid sha256:bd276b95419a1fd8f44a1e50dbf59f8229bd9212c44b9d081741c8302607df38
size 7288
