version https://git-lfs.github.com/spec/v1
oid sha256:7d0aa3682de9e1e743ece0f718502daadd3c3740f85723e2c3be7c19f7e357d5
size 6136
