version https://git-lfs.github.com/spec/v1
oid sha256:76c1af31a10b216306d37ec30eb94395dcdf46f30429822dd907f47469ca4aad
size 43402
