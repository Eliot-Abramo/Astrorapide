version https://git-lfs.github.com/spec/v1
oid sha256:d9fd3eaf83db58d07ad955b81006a356376a587f56ba65c4e3a56e804b0c9a26
size 14328
