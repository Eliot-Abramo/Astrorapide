version https://git-lfs.github.com/spec/v1
oid sha256:a2392877b3b3763da9426d75f6c5ae6a69ffd68bbc1e04f77d27a6ade87a91b4
size 54842
