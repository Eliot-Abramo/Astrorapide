version https://git-lfs.github.com/spec/v1
oid sha256:7fa635bcc5f0178d971b2fed35ccf91de2e496318a64dadb5875fd5c6171ddb8
size 2107
