version https://git-lfs.github.com/spec/v1
oid sha256:1a21d32d9880fd78360c3c0358f921d0c54e24003e058fa071255fc46fe8f29e
size 24272
