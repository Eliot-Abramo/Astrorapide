version https://git-lfs.github.com/spec/v1
oid sha256:a9feffb6494273b63936912baf61bb510ee68ad26169a7ac9fa980d875d39544
size 1508
