version https://git-lfs.github.com/spec/v1
oid sha256:243a279b7e44962e361c9e4dc91fee1ab0fe88a3f02b96c8b817acc8862835c5
size 2103
