version https://git-lfs.github.com/spec/v1
oid sha256:c956445108ef983142e9191288c0e5b3831cc3b9aa16fcb47bb0449c4fb24100
size 39044
