version https://git-lfs.github.com/spec/v1
oid sha256:40e719de4a2103a09b0dbc3e4a005438026d9fc79fba941566d0245c657ac2f9
size 14489
