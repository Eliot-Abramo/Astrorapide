version https://git-lfs.github.com/spec/v1
oid sha256:ba0d61831946f3246ac3fdddc34bca963564810b4a1dc8d8e5c141e63966310e
size 4477
