version https://git-lfs.github.com/spec/v1
oid sha256:c6c221dac68ddf48b93b32aa94b22cd8cf007ee5f916ab089b3aee2a7261a7b0
size 2107
