version https://git-lfs.github.com/spec/v1
oid sha256:7c3930050f34a4922fb270dc229a9689f8967d25fd98adce0772794767b9312b
size 54937
