version https://git-lfs.github.com/spec/v1
oid sha256:a822644279f877998803e2c019c40c4c2eb76c3607a609234452cf485fbf10bf
size 38790
