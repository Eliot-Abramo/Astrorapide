version https://git-lfs.github.com/spec/v1
oid sha256:29dd2de4869fc331c72353b4ef8d7e031c1c227651cc52847bd6d9d960627a78
size 44499
