version https://git-lfs.github.com/spec/v1
oid sha256:708d60fa131866e90536ee6fe0fe94742d06593b5033c21d02f41bd3c4665469
size 1508
