version https://git-lfs.github.com/spec/v1
oid sha256:dc7487c36854171873e2771536ceed48c618f9dcf43bc9e305d0fcb93d7caace
size 5345
