version https://git-lfs.github.com/spec/v1
oid sha256:2481ca71a8b70ea47037124065ff37ada0f1d066f7cef884eabf1f4ad5c75527
size 13401
