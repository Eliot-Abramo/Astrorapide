version https://git-lfs.github.com/spec/v1
oid sha256:91c0726e7f2f8eaafc6158f832de08e8eba71a24e336697f24cbe8f3244f2003
size 2116
