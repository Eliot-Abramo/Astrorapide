version https://git-lfs.github.com/spec/v1
oid sha256:d498b0eec913bbf8812335584c21ea45637b128029fe568de1f9f2220cec1319
size 3989
