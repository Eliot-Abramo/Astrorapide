version https://git-lfs.github.com/spec/v1
oid sha256:b0cd1d968c8dbd4a47b46b4c2a94c4185da645bb862c3c2e409da268bb96182e
size 2836
