version https://git-lfs.github.com/spec/v1
oid sha256:a3291968729f9fc0fa423d85c54077f063ea36ef5fbf4cbda34e481d028e6ca5
size 19571
