version https://git-lfs.github.com/spec/v1
oid sha256:542146892f61b644e143c8133dc21c213cba5483c261b8df1e075792d125c151
size 47638
