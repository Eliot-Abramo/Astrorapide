version https://git-lfs.github.com/spec/v1
oid sha256:fe7e96d7588a2e9549be752b9ed1abb05eb6dd474aed17696098539d2aaa8b24
size 51998
