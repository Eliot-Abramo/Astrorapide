version https://git-lfs.github.com/spec/v1
oid sha256:87c40caea7665de79f1213ad0cfc1be574609a71f2f6d84e5ceb02e60f8b8de6
size 2851
