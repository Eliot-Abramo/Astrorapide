version https://git-lfs.github.com/spec/v1
oid sha256:f3c65274720b602d45b7e362ac95439f8cf4365555a968e5e92a6c24cacf98e6
size 43936
