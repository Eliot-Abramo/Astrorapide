version https://git-lfs.github.com/spec/v1
oid sha256:c39f738bf89f7dacf649e4e3164258a535a0826e8f3fffb8a9ae857de73e27c9
size 13484
