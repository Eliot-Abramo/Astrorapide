version https://git-lfs.github.com/spec/v1
oid sha256:d6c8c86644ef0ccd1fceff0ba850547c56348027450db5eaf954c4dc6c7760c2
size 14417
