version https://git-lfs.github.com/spec/v1
oid sha256:2e6142a668db437f4fe0a75b7559151c2b28a140c2e66caec5e32d156898a451
size 3619
