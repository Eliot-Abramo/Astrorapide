version https://git-lfs.github.com/spec/v1
oid sha256:96e1e8e77ef7bf7da41359b9f49210c44e2cbf42a96d274fd28b7806b63b4952
size 1823
