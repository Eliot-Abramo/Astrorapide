version https://git-lfs.github.com/spec/v1
oid sha256:6903e47687b2c8b532835f9b2d6f845c3fa4b0bae0653c4424c714645cd8a989
size 43954
