version https://git-lfs.github.com/spec/v1
oid sha256:d8dff8901f8e623faa65f2065768cc03fb3d46d099b505d9c980218435ca2c11
size 2420
