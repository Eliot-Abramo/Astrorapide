version https://git-lfs.github.com/spec/v1
oid sha256:530b585b022320db8ddcc8aebdb93e29b0ef3a742f0c553e1449a9004a1e4b7c
size 7284
