version https://git-lfs.github.com/spec/v1
oid sha256:08d661077584f1bd6c19e1f2dfe6c326a5f25c74a368a7ec137cdc1aad9c1679
size 16968
