version https://git-lfs.github.com/spec/v1
oid sha256:0b66c4c679fbb8615c6a117d353ae657f25ca85783b86a3e0cd5077b6ab7a781
size 1867
