version https://git-lfs.github.com/spec/v1
oid sha256:41fe58cefe1d154327db65acd22c262bb2f002586c82447fdc3daf6bb9dce063
size 1817
