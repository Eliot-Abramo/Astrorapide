version https://git-lfs.github.com/spec/v1
oid sha256:59fccc684a7fbbed9e86ebda928fa7ea2d7b86800487a0151d310f8447fffa79
size 2844
