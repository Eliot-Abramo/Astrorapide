version https://git-lfs.github.com/spec/v1
oid sha256:4591eba3446401b1df1c246fedb45eeb14ad1cad01b28356f7aeb10fd15ed2f5
size 76095
