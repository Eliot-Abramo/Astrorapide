version https://git-lfs.github.com/spec/v1
oid sha256:dafc6cea6299adaccc30c03324671a7fb21189ac0198c22b4beef847bfa95176
size 2111
