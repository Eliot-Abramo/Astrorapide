version https://git-lfs.github.com/spec/v1
oid sha256:60483bdc2387c10eda01dd54cb7236f4339e0a05fb3479cfdb9fa61f034e4cdc
size 16975
