version https://git-lfs.github.com/spec/v1
oid sha256:c1b94f8b6e869ee6251c7e5c1f94094f394ed7acb85afea562e6ad0303e8af7c
size 13359
