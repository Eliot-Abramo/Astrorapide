version https://git-lfs.github.com/spec/v1
oid sha256:52df25698049d77b0e57ac99d3dc966b55c16d8090f458bf6564b004cafd48bc
size 2108
