version https://git-lfs.github.com/spec/v1
oid sha256:44fc0cac1f1b6079fc9db34abf3bd3f8189cdce5a314813aed7d76a83774494a
size 14486
