version https://git-lfs.github.com/spec/v1
oid sha256:6e7ebe3606ba209f92b905737d221c29a1c57e14ab88df04cde65c5711935c5d
size 54937
