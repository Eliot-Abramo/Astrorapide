version https://git-lfs.github.com/spec/v1
oid sha256:88d1dbe62b1684b56740394d7b9517f93a230dffab01afba129ba775cff4f650
size 13365
