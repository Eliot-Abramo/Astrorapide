version https://git-lfs.github.com/spec/v1
oid sha256:d50e6cb18f7bea358a2c271f53c230a0a9dd77a8242816a8c058ee4de735ab6e
size 54769
