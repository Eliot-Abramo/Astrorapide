version https://git-lfs.github.com/spec/v1
oid sha256:56cdf8c4bc9626aefbefc4c1024e2781a7c864a7fb70b2d77a4844d175c83a84
size 60942
